 module MUL #(vparam1, vparam2, vparamN)(
 port1,
 port2,
 portN
 );
BASIC #(.vparamB1(19), .vparamB2(6), .vparamBN(5)) BASIC1 (.portBA1(xxx), .portBA2(yyy));
 start of module MUL
 middle of module MUL
 end of module MUL
 endmodule
