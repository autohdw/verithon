 module Delay0000000009 (
    i_data, o_data
 );
 // Input and output ports
 input [14-1:0] i_data;
 output [14-1:0] o_data;
 assign o_data = i_data;
 endmodule
