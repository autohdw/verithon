 module BASIC #(vparamB1, vparamB2, vparamBN)(
 portBA1,
 portBA2,
 );
 start of module BASIC
 middle of module BASIC
 end of module BASIC
 endmodule
