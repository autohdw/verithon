 module M2V0000000001 (
     i_matrix, i_vector, o_result,
     i_clk
 );
 input wire [2*256*4*12-1:0] i_matrix;
 input wire [2*4*12-1:0] i_vector;
 output wire [2*256*12-1:0] o_result;
 input wire i_clk;
 wire [256*4*12-1:0] matrix_r, matrix_i;
 wire [4*12-1:0] vector_r, vector_i;
 assign matrix_r = i_matrix[256*4*12-1:0];
 assign matrix_i = i_matrix[2*256*4*12-1:256*4*12];
 assign vector_r = i_vector[4*12-1:0];
 assign vector_i = i_vector[2*4*12-1:4*12];
 // Layer 1: Add and Sub
 wire [13-1:0] a_plus_b [0:4-1];
 wire [13-1:0] b_minus_a [0:4-1];
 wire [13-1:0] c_plus_d [0:256-1][0:4-1];
Add0000000001  u_0000000001_Add0000000001(.i_data_1(vector_r[0*12+:12]), .i_data_2(vector_i[0*12+:12]), .o_data(a_plus_b[0]), .i_clk(i_clk));
Sub0000000001  u_0000000001_Sub0000000001(.i_data_1(vector_i[0*12+:12]), .i_data_2(vector_r[0*12+:12]), .o_data(b_minus_a[0]), .i_clk(i_clk));
Add0000000001  u_0000000002_Add0000000001(.i_data_1(matrix_r[0*12+:12]), .i_data_2(matrix_i[0*12+:12]), .o_data(c_plus_d[0][0]), .i_clk(i_clk));
Add0000000001  u_0000000003_Add0000000001(.i_data_1(matrix_r[1*12+:12]), .i_data_2(matrix_i[1*12+:12]), .o_data(c_plus_d[1][0]), .i_clk(i_clk));
Add0000000001  u_0000000004_Add0000000001(.i_data_1(matrix_r[2*12+:12]), .i_data_2(matrix_i[2*12+:12]), .o_data(c_plus_d[2][0]), .i_clk(i_clk));
Add0000000001  u_0000000005_Add0000000001(.i_data_1(matrix_r[3*12+:12]), .i_data_2(matrix_i[3*12+:12]), .o_data(c_plus_d[3][0]), .i_clk(i_clk));
Add0000000001  u_0000000006_Add0000000001(.i_data_1(matrix_r[4*12+:12]), .i_data_2(matrix_i[4*12+:12]), .o_data(c_plus_d[4][0]), .i_clk(i_clk));
Add0000000001  u_0000000007_Add0000000001(.i_data_1(matrix_r[5*12+:12]), .i_data_2(matrix_i[5*12+:12]), .o_data(c_plus_d[5][0]), .i_clk(i_clk));
Add0000000001  u_0000000008_Add0000000001(.i_data_1(matrix_r[6*12+:12]), .i_data_2(matrix_i[6*12+:12]), .o_data(c_plus_d[6][0]), .i_clk(i_clk));
Add0000000001  u_0000000009_Add0000000001(.i_data_1(matrix_r[7*12+:12]), .i_data_2(matrix_i[7*12+:12]), .o_data(c_plus_d[7][0]), .i_clk(i_clk));
Add0000000001  u_000000000A_Add0000000001(.i_data_1(matrix_r[8*12+:12]), .i_data_2(matrix_i[8*12+:12]), .o_data(c_plus_d[8][0]), .i_clk(i_clk));
Add0000000001  u_000000000B_Add0000000001(.i_data_1(matrix_r[9*12+:12]), .i_data_2(matrix_i[9*12+:12]), .o_data(c_plus_d[9][0]), .i_clk(i_clk));
Add0000000001  u_000000000C_Add0000000001(.i_data_1(matrix_r[10*12+:12]), .i_data_2(matrix_i[10*12+:12]), .o_data(c_plus_d[10][0]), .i_clk(i_clk));
Add0000000001  u_000000000D_Add0000000001(.i_data_1(matrix_r[11*12+:12]), .i_data_2(matrix_i[11*12+:12]), .o_data(c_plus_d[11][0]), .i_clk(i_clk));
Add0000000001  u_000000000E_Add0000000001(.i_data_1(matrix_r[12*12+:12]), .i_data_2(matrix_i[12*12+:12]), .o_data(c_plus_d[12][0]), .i_clk(i_clk));
Add0000000001  u_000000000F_Add0000000001(.i_data_1(matrix_r[13*12+:12]), .i_data_2(matrix_i[13*12+:12]), .o_data(c_plus_d[13][0]), .i_clk(i_clk));
Add0000000001  u_0000000010_Add0000000001(.i_data_1(matrix_r[14*12+:12]), .i_data_2(matrix_i[14*12+:12]), .o_data(c_plus_d[14][0]), .i_clk(i_clk));
Add0000000001  u_0000000011_Add0000000001(.i_data_1(matrix_r[15*12+:12]), .i_data_2(matrix_i[15*12+:12]), .o_data(c_plus_d[15][0]), .i_clk(i_clk));
Add0000000001  u_0000000012_Add0000000001(.i_data_1(matrix_r[16*12+:12]), .i_data_2(matrix_i[16*12+:12]), .o_data(c_plus_d[16][0]), .i_clk(i_clk));
Add0000000001  u_0000000013_Add0000000001(.i_data_1(matrix_r[17*12+:12]), .i_data_2(matrix_i[17*12+:12]), .o_data(c_plus_d[17][0]), .i_clk(i_clk));
Add0000000001  u_0000000014_Add0000000001(.i_data_1(matrix_r[18*12+:12]), .i_data_2(matrix_i[18*12+:12]), .o_data(c_plus_d[18][0]), .i_clk(i_clk));
Add0000000001  u_0000000015_Add0000000001(.i_data_1(matrix_r[19*12+:12]), .i_data_2(matrix_i[19*12+:12]), .o_data(c_plus_d[19][0]), .i_clk(i_clk));
Add0000000001  u_0000000016_Add0000000001(.i_data_1(matrix_r[20*12+:12]), .i_data_2(matrix_i[20*12+:12]), .o_data(c_plus_d[20][0]), .i_clk(i_clk));
Add0000000001  u_0000000017_Add0000000001(.i_data_1(matrix_r[21*12+:12]), .i_data_2(matrix_i[21*12+:12]), .o_data(c_plus_d[21][0]), .i_clk(i_clk));
Add0000000001  u_0000000018_Add0000000001(.i_data_1(matrix_r[22*12+:12]), .i_data_2(matrix_i[22*12+:12]), .o_data(c_plus_d[22][0]), .i_clk(i_clk));
Add0000000001  u_0000000019_Add0000000001(.i_data_1(matrix_r[23*12+:12]), .i_data_2(matrix_i[23*12+:12]), .o_data(c_plus_d[23][0]), .i_clk(i_clk));
Add0000000001  u_000000001A_Add0000000001(.i_data_1(matrix_r[24*12+:12]), .i_data_2(matrix_i[24*12+:12]), .o_data(c_plus_d[24][0]), .i_clk(i_clk));
Add0000000001  u_000000001B_Add0000000001(.i_data_1(matrix_r[25*12+:12]), .i_data_2(matrix_i[25*12+:12]), .o_data(c_plus_d[25][0]), .i_clk(i_clk));
Add0000000001  u_000000001C_Add0000000001(.i_data_1(matrix_r[26*12+:12]), .i_data_2(matrix_i[26*12+:12]), .o_data(c_plus_d[26][0]), .i_clk(i_clk));
Add0000000001  u_000000001D_Add0000000001(.i_data_1(matrix_r[27*12+:12]), .i_data_2(matrix_i[27*12+:12]), .o_data(c_plus_d[27][0]), .i_clk(i_clk));
Add0000000001  u_000000001E_Add0000000001(.i_data_1(matrix_r[28*12+:12]), .i_data_2(matrix_i[28*12+:12]), .o_data(c_plus_d[28][0]), .i_clk(i_clk));
Add0000000001  u_000000001F_Add0000000001(.i_data_1(matrix_r[29*12+:12]), .i_data_2(matrix_i[29*12+:12]), .o_data(c_plus_d[29][0]), .i_clk(i_clk));
Add0000000001  u_0000000020_Add0000000001(.i_data_1(matrix_r[30*12+:12]), .i_data_2(matrix_i[30*12+:12]), .o_data(c_plus_d[30][0]), .i_clk(i_clk));
Add0000000001  u_0000000021_Add0000000001(.i_data_1(matrix_r[31*12+:12]), .i_data_2(matrix_i[31*12+:12]), .o_data(c_plus_d[31][0]), .i_clk(i_clk));
Add0000000001  u_0000000022_Add0000000001(.i_data_1(matrix_r[32*12+:12]), .i_data_2(matrix_i[32*12+:12]), .o_data(c_plus_d[32][0]), .i_clk(i_clk));
Add0000000001  u_0000000023_Add0000000001(.i_data_1(matrix_r[33*12+:12]), .i_data_2(matrix_i[33*12+:12]), .o_data(c_plus_d[33][0]), .i_clk(i_clk));
Add0000000001  u_0000000024_Add0000000001(.i_data_1(matrix_r[34*12+:12]), .i_data_2(matrix_i[34*12+:12]), .o_data(c_plus_d[34][0]), .i_clk(i_clk));
Add0000000001  u_0000000025_Add0000000001(.i_data_1(matrix_r[35*12+:12]), .i_data_2(matrix_i[35*12+:12]), .o_data(c_plus_d[35][0]), .i_clk(i_clk));
Add0000000001  u_0000000026_Add0000000001(.i_data_1(matrix_r[36*12+:12]), .i_data_2(matrix_i[36*12+:12]), .o_data(c_plus_d[36][0]), .i_clk(i_clk));
Add0000000001  u_0000000027_Add0000000001(.i_data_1(matrix_r[37*12+:12]), .i_data_2(matrix_i[37*12+:12]), .o_data(c_plus_d[37][0]), .i_clk(i_clk));
Add0000000001  u_0000000028_Add0000000001(.i_data_1(matrix_r[38*12+:12]), .i_data_2(matrix_i[38*12+:12]), .o_data(c_plus_d[38][0]), .i_clk(i_clk));
Add0000000001  u_0000000029_Add0000000001(.i_data_1(matrix_r[39*12+:12]), .i_data_2(matrix_i[39*12+:12]), .o_data(c_plus_d[39][0]), .i_clk(i_clk));
Add0000000001  u_000000002A_Add0000000001(.i_data_1(matrix_r[40*12+:12]), .i_data_2(matrix_i[40*12+:12]), .o_data(c_plus_d[40][0]), .i_clk(i_clk));
Add0000000001  u_000000002B_Add0000000001(.i_data_1(matrix_r[41*12+:12]), .i_data_2(matrix_i[41*12+:12]), .o_data(c_plus_d[41][0]), .i_clk(i_clk));
Add0000000001  u_000000002C_Add0000000001(.i_data_1(matrix_r[42*12+:12]), .i_data_2(matrix_i[42*12+:12]), .o_data(c_plus_d[42][0]), .i_clk(i_clk));
Add0000000001  u_000000002D_Add0000000001(.i_data_1(matrix_r[43*12+:12]), .i_data_2(matrix_i[43*12+:12]), .o_data(c_plus_d[43][0]), .i_clk(i_clk));
Add0000000001  u_000000002E_Add0000000001(.i_data_1(matrix_r[44*12+:12]), .i_data_2(matrix_i[44*12+:12]), .o_data(c_plus_d[44][0]), .i_clk(i_clk));
Add0000000001  u_000000002F_Add0000000001(.i_data_1(matrix_r[45*12+:12]), .i_data_2(matrix_i[45*12+:12]), .o_data(c_plus_d[45][0]), .i_clk(i_clk));
Add0000000001  u_0000000030_Add0000000001(.i_data_1(matrix_r[46*12+:12]), .i_data_2(matrix_i[46*12+:12]), .o_data(c_plus_d[46][0]), .i_clk(i_clk));
Add0000000001  u_0000000031_Add0000000001(.i_data_1(matrix_r[47*12+:12]), .i_data_2(matrix_i[47*12+:12]), .o_data(c_plus_d[47][0]), .i_clk(i_clk));
Add0000000001  u_0000000032_Add0000000001(.i_data_1(matrix_r[48*12+:12]), .i_data_2(matrix_i[48*12+:12]), .o_data(c_plus_d[48][0]), .i_clk(i_clk));
Add0000000001  u_0000000033_Add0000000001(.i_data_1(matrix_r[49*12+:12]), .i_data_2(matrix_i[49*12+:12]), .o_data(c_plus_d[49][0]), .i_clk(i_clk));
Add0000000001  u_0000000034_Add0000000001(.i_data_1(matrix_r[50*12+:12]), .i_data_2(matrix_i[50*12+:12]), .o_data(c_plus_d[50][0]), .i_clk(i_clk));
Add0000000001  u_0000000035_Add0000000001(.i_data_1(matrix_r[51*12+:12]), .i_data_2(matrix_i[51*12+:12]), .o_data(c_plus_d[51][0]), .i_clk(i_clk));
Add0000000001  u_0000000036_Add0000000001(.i_data_1(matrix_r[52*12+:12]), .i_data_2(matrix_i[52*12+:12]), .o_data(c_plus_d[52][0]), .i_clk(i_clk));
Add0000000001  u_0000000037_Add0000000001(.i_data_1(matrix_r[53*12+:12]), .i_data_2(matrix_i[53*12+:12]), .o_data(c_plus_d[53][0]), .i_clk(i_clk));
Add0000000001  u_0000000038_Add0000000001(.i_data_1(matrix_r[54*12+:12]), .i_data_2(matrix_i[54*12+:12]), .o_data(c_plus_d[54][0]), .i_clk(i_clk));
Add0000000001  u_0000000039_Add0000000001(.i_data_1(matrix_r[55*12+:12]), .i_data_2(matrix_i[55*12+:12]), .o_data(c_plus_d[55][0]), .i_clk(i_clk));
Add0000000001  u_000000003A_Add0000000001(.i_data_1(matrix_r[56*12+:12]), .i_data_2(matrix_i[56*12+:12]), .o_data(c_plus_d[56][0]), .i_clk(i_clk));
Add0000000001  u_000000003B_Add0000000001(.i_data_1(matrix_r[57*12+:12]), .i_data_2(matrix_i[57*12+:12]), .o_data(c_plus_d[57][0]), .i_clk(i_clk));
Add0000000001  u_000000003C_Add0000000001(.i_data_1(matrix_r[58*12+:12]), .i_data_2(matrix_i[58*12+:12]), .o_data(c_plus_d[58][0]), .i_clk(i_clk));
Add0000000001  u_000000003D_Add0000000001(.i_data_1(matrix_r[59*12+:12]), .i_data_2(matrix_i[59*12+:12]), .o_data(c_plus_d[59][0]), .i_clk(i_clk));
Add0000000001  u_000000003E_Add0000000001(.i_data_1(matrix_r[60*12+:12]), .i_data_2(matrix_i[60*12+:12]), .o_data(c_plus_d[60][0]), .i_clk(i_clk));
Add0000000001  u_000000003F_Add0000000001(.i_data_1(matrix_r[61*12+:12]), .i_data_2(matrix_i[61*12+:12]), .o_data(c_plus_d[61][0]), .i_clk(i_clk));
Add0000000001  u_0000000040_Add0000000001(.i_data_1(matrix_r[62*12+:12]), .i_data_2(matrix_i[62*12+:12]), .o_data(c_plus_d[62][0]), .i_clk(i_clk));
Add0000000001  u_0000000041_Add0000000001(.i_data_1(matrix_r[63*12+:12]), .i_data_2(matrix_i[63*12+:12]), .o_data(c_plus_d[63][0]), .i_clk(i_clk));
Add0000000001  u_0000000042_Add0000000001(.i_data_1(matrix_r[64*12+:12]), .i_data_2(matrix_i[64*12+:12]), .o_data(c_plus_d[64][0]), .i_clk(i_clk));
Add0000000001  u_0000000043_Add0000000001(.i_data_1(matrix_r[65*12+:12]), .i_data_2(matrix_i[65*12+:12]), .o_data(c_plus_d[65][0]), .i_clk(i_clk));
Add0000000001  u_0000000044_Add0000000001(.i_data_1(matrix_r[66*12+:12]), .i_data_2(matrix_i[66*12+:12]), .o_data(c_plus_d[66][0]), .i_clk(i_clk));
Add0000000001  u_0000000045_Add0000000001(.i_data_1(matrix_r[67*12+:12]), .i_data_2(matrix_i[67*12+:12]), .o_data(c_plus_d[67][0]), .i_clk(i_clk));
Add0000000001  u_0000000046_Add0000000001(.i_data_1(matrix_r[68*12+:12]), .i_data_2(matrix_i[68*12+:12]), .o_data(c_plus_d[68][0]), .i_clk(i_clk));
Add0000000001  u_0000000047_Add0000000001(.i_data_1(matrix_r[69*12+:12]), .i_data_2(matrix_i[69*12+:12]), .o_data(c_plus_d[69][0]), .i_clk(i_clk));
Add0000000001  u_0000000048_Add0000000001(.i_data_1(matrix_r[70*12+:12]), .i_data_2(matrix_i[70*12+:12]), .o_data(c_plus_d[70][0]), .i_clk(i_clk));
Add0000000001  u_0000000049_Add0000000001(.i_data_1(matrix_r[71*12+:12]), .i_data_2(matrix_i[71*12+:12]), .o_data(c_plus_d[71][0]), .i_clk(i_clk));
Add0000000001  u_000000004A_Add0000000001(.i_data_1(matrix_r[72*12+:12]), .i_data_2(matrix_i[72*12+:12]), .o_data(c_plus_d[72][0]), .i_clk(i_clk));
Add0000000001  u_000000004B_Add0000000001(.i_data_1(matrix_r[73*12+:12]), .i_data_2(matrix_i[73*12+:12]), .o_data(c_plus_d[73][0]), .i_clk(i_clk));
Add0000000001  u_000000004C_Add0000000001(.i_data_1(matrix_r[74*12+:12]), .i_data_2(matrix_i[74*12+:12]), .o_data(c_plus_d[74][0]), .i_clk(i_clk));
Add0000000001  u_000000004D_Add0000000001(.i_data_1(matrix_r[75*12+:12]), .i_data_2(matrix_i[75*12+:12]), .o_data(c_plus_d[75][0]), .i_clk(i_clk));
Add0000000001  u_000000004E_Add0000000001(.i_data_1(matrix_r[76*12+:12]), .i_data_2(matrix_i[76*12+:12]), .o_data(c_plus_d[76][0]), .i_clk(i_clk));
Add0000000001  u_000000004F_Add0000000001(.i_data_1(matrix_r[77*12+:12]), .i_data_2(matrix_i[77*12+:12]), .o_data(c_plus_d[77][0]), .i_clk(i_clk));
Add0000000001  u_0000000050_Add0000000001(.i_data_1(matrix_r[78*12+:12]), .i_data_2(matrix_i[78*12+:12]), .o_data(c_plus_d[78][0]), .i_clk(i_clk));
Add0000000001  u_0000000051_Add0000000001(.i_data_1(matrix_r[79*12+:12]), .i_data_2(matrix_i[79*12+:12]), .o_data(c_plus_d[79][0]), .i_clk(i_clk));
Add0000000001  u_0000000052_Add0000000001(.i_data_1(matrix_r[80*12+:12]), .i_data_2(matrix_i[80*12+:12]), .o_data(c_plus_d[80][0]), .i_clk(i_clk));
Add0000000001  u_0000000053_Add0000000001(.i_data_1(matrix_r[81*12+:12]), .i_data_2(matrix_i[81*12+:12]), .o_data(c_plus_d[81][0]), .i_clk(i_clk));
Add0000000001  u_0000000054_Add0000000001(.i_data_1(matrix_r[82*12+:12]), .i_data_2(matrix_i[82*12+:12]), .o_data(c_plus_d[82][0]), .i_clk(i_clk));
Add0000000001  u_0000000055_Add0000000001(.i_data_1(matrix_r[83*12+:12]), .i_data_2(matrix_i[83*12+:12]), .o_data(c_plus_d[83][0]), .i_clk(i_clk));
Add0000000001  u_0000000056_Add0000000001(.i_data_1(matrix_r[84*12+:12]), .i_data_2(matrix_i[84*12+:12]), .o_data(c_plus_d[84][0]), .i_clk(i_clk));
Add0000000001  u_0000000057_Add0000000001(.i_data_1(matrix_r[85*12+:12]), .i_data_2(matrix_i[85*12+:12]), .o_data(c_plus_d[85][0]), .i_clk(i_clk));
Add0000000001  u_0000000058_Add0000000001(.i_data_1(matrix_r[86*12+:12]), .i_data_2(matrix_i[86*12+:12]), .o_data(c_plus_d[86][0]), .i_clk(i_clk));
Add0000000001  u_0000000059_Add0000000001(.i_data_1(matrix_r[87*12+:12]), .i_data_2(matrix_i[87*12+:12]), .o_data(c_plus_d[87][0]), .i_clk(i_clk));
Add0000000001  u_000000005A_Add0000000001(.i_data_1(matrix_r[88*12+:12]), .i_data_2(matrix_i[88*12+:12]), .o_data(c_plus_d[88][0]), .i_clk(i_clk));
Add0000000001  u_000000005B_Add0000000001(.i_data_1(matrix_r[89*12+:12]), .i_data_2(matrix_i[89*12+:12]), .o_data(c_plus_d[89][0]), .i_clk(i_clk));
Add0000000001  u_000000005C_Add0000000001(.i_data_1(matrix_r[90*12+:12]), .i_data_2(matrix_i[90*12+:12]), .o_data(c_plus_d[90][0]), .i_clk(i_clk));
Add0000000001  u_000000005D_Add0000000001(.i_data_1(matrix_r[91*12+:12]), .i_data_2(matrix_i[91*12+:12]), .o_data(c_plus_d[91][0]), .i_clk(i_clk));
Add0000000001  u_000000005E_Add0000000001(.i_data_1(matrix_r[92*12+:12]), .i_data_2(matrix_i[92*12+:12]), .o_data(c_plus_d[92][0]), .i_clk(i_clk));
Add0000000001  u_000000005F_Add0000000001(.i_data_1(matrix_r[93*12+:12]), .i_data_2(matrix_i[93*12+:12]), .o_data(c_plus_d[93][0]), .i_clk(i_clk));
Add0000000001  u_0000000060_Add0000000001(.i_data_1(matrix_r[94*12+:12]), .i_data_2(matrix_i[94*12+:12]), .o_data(c_plus_d[94][0]), .i_clk(i_clk));
Add0000000001  u_0000000061_Add0000000001(.i_data_1(matrix_r[95*12+:12]), .i_data_2(matrix_i[95*12+:12]), .o_data(c_plus_d[95][0]), .i_clk(i_clk));
Add0000000001  u_0000000062_Add0000000001(.i_data_1(matrix_r[96*12+:12]), .i_data_2(matrix_i[96*12+:12]), .o_data(c_plus_d[96][0]), .i_clk(i_clk));
Add0000000001  u_0000000063_Add0000000001(.i_data_1(matrix_r[97*12+:12]), .i_data_2(matrix_i[97*12+:12]), .o_data(c_plus_d[97][0]), .i_clk(i_clk));
Add0000000001  u_0000000064_Add0000000001(.i_data_1(matrix_r[98*12+:12]), .i_data_2(matrix_i[98*12+:12]), .o_data(c_plus_d[98][0]), .i_clk(i_clk));
Add0000000001  u_0000000065_Add0000000001(.i_data_1(matrix_r[99*12+:12]), .i_data_2(matrix_i[99*12+:12]), .o_data(c_plus_d[99][0]), .i_clk(i_clk));
Add0000000001  u_0000000066_Add0000000001(.i_data_1(matrix_r[100*12+:12]), .i_data_2(matrix_i[100*12+:12]), .o_data(c_plus_d[100][0]), .i_clk(i_clk));
Add0000000001  u_0000000067_Add0000000001(.i_data_1(matrix_r[101*12+:12]), .i_data_2(matrix_i[101*12+:12]), .o_data(c_plus_d[101][0]), .i_clk(i_clk));
Add0000000001  u_0000000068_Add0000000001(.i_data_1(matrix_r[102*12+:12]), .i_data_2(matrix_i[102*12+:12]), .o_data(c_plus_d[102][0]), .i_clk(i_clk));
Add0000000001  u_0000000069_Add0000000001(.i_data_1(matrix_r[103*12+:12]), .i_data_2(matrix_i[103*12+:12]), .o_data(c_plus_d[103][0]), .i_clk(i_clk));
Add0000000001  u_000000006A_Add0000000001(.i_data_1(matrix_r[104*12+:12]), .i_data_2(matrix_i[104*12+:12]), .o_data(c_plus_d[104][0]), .i_clk(i_clk));
Add0000000001  u_000000006B_Add0000000001(.i_data_1(matrix_r[105*12+:12]), .i_data_2(matrix_i[105*12+:12]), .o_data(c_plus_d[105][0]), .i_clk(i_clk));
Add0000000001  u_000000006C_Add0000000001(.i_data_1(matrix_r[106*12+:12]), .i_data_2(matrix_i[106*12+:12]), .o_data(c_plus_d[106][0]), .i_clk(i_clk));
Add0000000001  u_000000006D_Add0000000001(.i_data_1(matrix_r[107*12+:12]), .i_data_2(matrix_i[107*12+:12]), .o_data(c_plus_d[107][0]), .i_clk(i_clk));
Add0000000001  u_000000006E_Add0000000001(.i_data_1(matrix_r[108*12+:12]), .i_data_2(matrix_i[108*12+:12]), .o_data(c_plus_d[108][0]), .i_clk(i_clk));
Add0000000001  u_000000006F_Add0000000001(.i_data_1(matrix_r[109*12+:12]), .i_data_2(matrix_i[109*12+:12]), .o_data(c_plus_d[109][0]), .i_clk(i_clk));
Add0000000001  u_0000000070_Add0000000001(.i_data_1(matrix_r[110*12+:12]), .i_data_2(matrix_i[110*12+:12]), .o_data(c_plus_d[110][0]), .i_clk(i_clk));
Add0000000001  u_0000000071_Add0000000001(.i_data_1(matrix_r[111*12+:12]), .i_data_2(matrix_i[111*12+:12]), .o_data(c_plus_d[111][0]), .i_clk(i_clk));
Add0000000001  u_0000000072_Add0000000001(.i_data_1(matrix_r[112*12+:12]), .i_data_2(matrix_i[112*12+:12]), .o_data(c_plus_d[112][0]), .i_clk(i_clk));
Add0000000001  u_0000000073_Add0000000001(.i_data_1(matrix_r[113*12+:12]), .i_data_2(matrix_i[113*12+:12]), .o_data(c_plus_d[113][0]), .i_clk(i_clk));
Add0000000001  u_0000000074_Add0000000001(.i_data_1(matrix_r[114*12+:12]), .i_data_2(matrix_i[114*12+:12]), .o_data(c_plus_d[114][0]), .i_clk(i_clk));
Add0000000001  u_0000000075_Add0000000001(.i_data_1(matrix_r[115*12+:12]), .i_data_2(matrix_i[115*12+:12]), .o_data(c_plus_d[115][0]), .i_clk(i_clk));
Add0000000001  u_0000000076_Add0000000001(.i_data_1(matrix_r[116*12+:12]), .i_data_2(matrix_i[116*12+:12]), .o_data(c_plus_d[116][0]), .i_clk(i_clk));
Add0000000001  u_0000000077_Add0000000001(.i_data_1(matrix_r[117*12+:12]), .i_data_2(matrix_i[117*12+:12]), .o_data(c_plus_d[117][0]), .i_clk(i_clk));
Add0000000001  u_0000000078_Add0000000001(.i_data_1(matrix_r[118*12+:12]), .i_data_2(matrix_i[118*12+:12]), .o_data(c_plus_d[118][0]), .i_clk(i_clk));
Add0000000001  u_0000000079_Add0000000001(.i_data_1(matrix_r[119*12+:12]), .i_data_2(matrix_i[119*12+:12]), .o_data(c_plus_d[119][0]), .i_clk(i_clk));
Add0000000001  u_000000007A_Add0000000001(.i_data_1(matrix_r[120*12+:12]), .i_data_2(matrix_i[120*12+:12]), .o_data(c_plus_d[120][0]), .i_clk(i_clk));
Add0000000001  u_000000007B_Add0000000001(.i_data_1(matrix_r[121*12+:12]), .i_data_2(matrix_i[121*12+:12]), .o_data(c_plus_d[121][0]), .i_clk(i_clk));
Add0000000001  u_000000007C_Add0000000001(.i_data_1(matrix_r[122*12+:12]), .i_data_2(matrix_i[122*12+:12]), .o_data(c_plus_d[122][0]), .i_clk(i_clk));
Add0000000001  u_000000007D_Add0000000001(.i_data_1(matrix_r[123*12+:12]), .i_data_2(matrix_i[123*12+:12]), .o_data(c_plus_d[123][0]), .i_clk(i_clk));
Add0000000001  u_000000007E_Add0000000001(.i_data_1(matrix_r[124*12+:12]), .i_data_2(matrix_i[124*12+:12]), .o_data(c_plus_d[124][0]), .i_clk(i_clk));
Add0000000001  u_000000007F_Add0000000001(.i_data_1(matrix_r[125*12+:12]), .i_data_2(matrix_i[125*12+:12]), .o_data(c_plus_d[125][0]), .i_clk(i_clk));
Add0000000001  u_0000000080_Add0000000001(.i_data_1(matrix_r[126*12+:12]), .i_data_2(matrix_i[126*12+:12]), .o_data(c_plus_d[126][0]), .i_clk(i_clk));
Add0000000001  u_0000000081_Add0000000001(.i_data_1(matrix_r[127*12+:12]), .i_data_2(matrix_i[127*12+:12]), .o_data(c_plus_d[127][0]), .i_clk(i_clk));
Add0000000001  u_0000000082_Add0000000001(.i_data_1(matrix_r[128*12+:12]), .i_data_2(matrix_i[128*12+:12]), .o_data(c_plus_d[128][0]), .i_clk(i_clk));
Add0000000001  u_0000000083_Add0000000001(.i_data_1(matrix_r[129*12+:12]), .i_data_2(matrix_i[129*12+:12]), .o_data(c_plus_d[129][0]), .i_clk(i_clk));
Add0000000001  u_0000000084_Add0000000001(.i_data_1(matrix_r[130*12+:12]), .i_data_2(matrix_i[130*12+:12]), .o_data(c_plus_d[130][0]), .i_clk(i_clk));
Add0000000001  u_0000000085_Add0000000001(.i_data_1(matrix_r[131*12+:12]), .i_data_2(matrix_i[131*12+:12]), .o_data(c_plus_d[131][0]), .i_clk(i_clk));
Add0000000001  u_0000000086_Add0000000001(.i_data_1(matrix_r[132*12+:12]), .i_data_2(matrix_i[132*12+:12]), .o_data(c_plus_d[132][0]), .i_clk(i_clk));
Add0000000001  u_0000000087_Add0000000001(.i_data_1(matrix_r[133*12+:12]), .i_data_2(matrix_i[133*12+:12]), .o_data(c_plus_d[133][0]), .i_clk(i_clk));
Add0000000001  u_0000000088_Add0000000001(.i_data_1(matrix_r[134*12+:12]), .i_data_2(matrix_i[134*12+:12]), .o_data(c_plus_d[134][0]), .i_clk(i_clk));
Add0000000001  u_0000000089_Add0000000001(.i_data_1(matrix_r[135*12+:12]), .i_data_2(matrix_i[135*12+:12]), .o_data(c_plus_d[135][0]), .i_clk(i_clk));
Add0000000001  u_000000008A_Add0000000001(.i_data_1(matrix_r[136*12+:12]), .i_data_2(matrix_i[136*12+:12]), .o_data(c_plus_d[136][0]), .i_clk(i_clk));
Add0000000001  u_000000008B_Add0000000001(.i_data_1(matrix_r[137*12+:12]), .i_data_2(matrix_i[137*12+:12]), .o_data(c_plus_d[137][0]), .i_clk(i_clk));
Add0000000001  u_000000008C_Add0000000001(.i_data_1(matrix_r[138*12+:12]), .i_data_2(matrix_i[138*12+:12]), .o_data(c_plus_d[138][0]), .i_clk(i_clk));
Add0000000001  u_000000008D_Add0000000001(.i_data_1(matrix_r[139*12+:12]), .i_data_2(matrix_i[139*12+:12]), .o_data(c_plus_d[139][0]), .i_clk(i_clk));
Add0000000001  u_000000008E_Add0000000001(.i_data_1(matrix_r[140*12+:12]), .i_data_2(matrix_i[140*12+:12]), .o_data(c_plus_d[140][0]), .i_clk(i_clk));
Add0000000001  u_000000008F_Add0000000001(.i_data_1(matrix_r[141*12+:12]), .i_data_2(matrix_i[141*12+:12]), .o_data(c_plus_d[141][0]), .i_clk(i_clk));
Add0000000001  u_0000000090_Add0000000001(.i_data_1(matrix_r[142*12+:12]), .i_data_2(matrix_i[142*12+:12]), .o_data(c_plus_d[142][0]), .i_clk(i_clk));
Add0000000001  u_0000000091_Add0000000001(.i_data_1(matrix_r[143*12+:12]), .i_data_2(matrix_i[143*12+:12]), .o_data(c_plus_d[143][0]), .i_clk(i_clk));
Add0000000001  u_0000000092_Add0000000001(.i_data_1(matrix_r[144*12+:12]), .i_data_2(matrix_i[144*12+:12]), .o_data(c_plus_d[144][0]), .i_clk(i_clk));
Add0000000001  u_0000000093_Add0000000001(.i_data_1(matrix_r[145*12+:12]), .i_data_2(matrix_i[145*12+:12]), .o_data(c_plus_d[145][0]), .i_clk(i_clk));
Add0000000001  u_0000000094_Add0000000001(.i_data_1(matrix_r[146*12+:12]), .i_data_2(matrix_i[146*12+:12]), .o_data(c_plus_d[146][0]), .i_clk(i_clk));
Add0000000001  u_0000000095_Add0000000001(.i_data_1(matrix_r[147*12+:12]), .i_data_2(matrix_i[147*12+:12]), .o_data(c_plus_d[147][0]), .i_clk(i_clk));
Add0000000001  u_0000000096_Add0000000001(.i_data_1(matrix_r[148*12+:12]), .i_data_2(matrix_i[148*12+:12]), .o_data(c_plus_d[148][0]), .i_clk(i_clk));
Add0000000001  u_0000000097_Add0000000001(.i_data_1(matrix_r[149*12+:12]), .i_data_2(matrix_i[149*12+:12]), .o_data(c_plus_d[149][0]), .i_clk(i_clk));
Add0000000001  u_0000000098_Add0000000001(.i_data_1(matrix_r[150*12+:12]), .i_data_2(matrix_i[150*12+:12]), .o_data(c_plus_d[150][0]), .i_clk(i_clk));
Add0000000001  u_0000000099_Add0000000001(.i_data_1(matrix_r[151*12+:12]), .i_data_2(matrix_i[151*12+:12]), .o_data(c_plus_d[151][0]), .i_clk(i_clk));
Add0000000001  u_000000009A_Add0000000001(.i_data_1(matrix_r[152*12+:12]), .i_data_2(matrix_i[152*12+:12]), .o_data(c_plus_d[152][0]), .i_clk(i_clk));
Add0000000001  u_000000009B_Add0000000001(.i_data_1(matrix_r[153*12+:12]), .i_data_2(matrix_i[153*12+:12]), .o_data(c_plus_d[153][0]), .i_clk(i_clk));
Add0000000001  u_000000009C_Add0000000001(.i_data_1(matrix_r[154*12+:12]), .i_data_2(matrix_i[154*12+:12]), .o_data(c_plus_d[154][0]), .i_clk(i_clk));
Add0000000001  u_000000009D_Add0000000001(.i_data_1(matrix_r[155*12+:12]), .i_data_2(matrix_i[155*12+:12]), .o_data(c_plus_d[155][0]), .i_clk(i_clk));
Add0000000001  u_000000009E_Add0000000001(.i_data_1(matrix_r[156*12+:12]), .i_data_2(matrix_i[156*12+:12]), .o_data(c_plus_d[156][0]), .i_clk(i_clk));
Add0000000001  u_000000009F_Add0000000001(.i_data_1(matrix_r[157*12+:12]), .i_data_2(matrix_i[157*12+:12]), .o_data(c_plus_d[157][0]), .i_clk(i_clk));
Add0000000001  u_00000000A0_Add0000000001(.i_data_1(matrix_r[158*12+:12]), .i_data_2(matrix_i[158*12+:12]), .o_data(c_plus_d[158][0]), .i_clk(i_clk));
Add0000000001  u_00000000A1_Add0000000001(.i_data_1(matrix_r[159*12+:12]), .i_data_2(matrix_i[159*12+:12]), .o_data(c_plus_d[159][0]), .i_clk(i_clk));
Add0000000001  u_00000000A2_Add0000000001(.i_data_1(matrix_r[160*12+:12]), .i_data_2(matrix_i[160*12+:12]), .o_data(c_plus_d[160][0]), .i_clk(i_clk));
Add0000000001  u_00000000A3_Add0000000001(.i_data_1(matrix_r[161*12+:12]), .i_data_2(matrix_i[161*12+:12]), .o_data(c_plus_d[161][0]), .i_clk(i_clk));
Add0000000001  u_00000000A4_Add0000000001(.i_data_1(matrix_r[162*12+:12]), .i_data_2(matrix_i[162*12+:12]), .o_data(c_plus_d[162][0]), .i_clk(i_clk));
Add0000000001  u_00000000A5_Add0000000001(.i_data_1(matrix_r[163*12+:12]), .i_data_2(matrix_i[163*12+:12]), .o_data(c_plus_d[163][0]), .i_clk(i_clk));
Add0000000001  u_00000000A6_Add0000000001(.i_data_1(matrix_r[164*12+:12]), .i_data_2(matrix_i[164*12+:12]), .o_data(c_plus_d[164][0]), .i_clk(i_clk));
Add0000000001  u_00000000A7_Add0000000001(.i_data_1(matrix_r[165*12+:12]), .i_data_2(matrix_i[165*12+:12]), .o_data(c_plus_d[165][0]), .i_clk(i_clk));
Add0000000001  u_00000000A8_Add0000000001(.i_data_1(matrix_r[166*12+:12]), .i_data_2(matrix_i[166*12+:12]), .o_data(c_plus_d[166][0]), .i_clk(i_clk));
Add0000000001  u_00000000A9_Add0000000001(.i_data_1(matrix_r[167*12+:12]), .i_data_2(matrix_i[167*12+:12]), .o_data(c_plus_d[167][0]), .i_clk(i_clk));
Add0000000001  u_00000000AA_Add0000000001(.i_data_1(matrix_r[168*12+:12]), .i_data_2(matrix_i[168*12+:12]), .o_data(c_plus_d[168][0]), .i_clk(i_clk));
Add0000000001  u_00000000AB_Add0000000001(.i_data_1(matrix_r[169*12+:12]), .i_data_2(matrix_i[169*12+:12]), .o_data(c_plus_d[169][0]), .i_clk(i_clk));
Add0000000001  u_00000000AC_Add0000000001(.i_data_1(matrix_r[170*12+:12]), .i_data_2(matrix_i[170*12+:12]), .o_data(c_plus_d[170][0]), .i_clk(i_clk));
Add0000000001  u_00000000AD_Add0000000001(.i_data_1(matrix_r[171*12+:12]), .i_data_2(matrix_i[171*12+:12]), .o_data(c_plus_d[171][0]), .i_clk(i_clk));
Add0000000001  u_00000000AE_Add0000000001(.i_data_1(matrix_r[172*12+:12]), .i_data_2(matrix_i[172*12+:12]), .o_data(c_plus_d[172][0]), .i_clk(i_clk));
Add0000000001  u_00000000AF_Add0000000001(.i_data_1(matrix_r[173*12+:12]), .i_data_2(matrix_i[173*12+:12]), .o_data(c_plus_d[173][0]), .i_clk(i_clk));
Add0000000001  u_00000000B0_Add0000000001(.i_data_1(matrix_r[174*12+:12]), .i_data_2(matrix_i[174*12+:12]), .o_data(c_plus_d[174][0]), .i_clk(i_clk));
Add0000000001  u_00000000B1_Add0000000001(.i_data_1(matrix_r[175*12+:12]), .i_data_2(matrix_i[175*12+:12]), .o_data(c_plus_d[175][0]), .i_clk(i_clk));
Add0000000001  u_00000000B2_Add0000000001(.i_data_1(matrix_r[176*12+:12]), .i_data_2(matrix_i[176*12+:12]), .o_data(c_plus_d[176][0]), .i_clk(i_clk));
Add0000000001  u_00000000B3_Add0000000001(.i_data_1(matrix_r[177*12+:12]), .i_data_2(matrix_i[177*12+:12]), .o_data(c_plus_d[177][0]), .i_clk(i_clk));
Add0000000001  u_00000000B4_Add0000000001(.i_data_1(matrix_r[178*12+:12]), .i_data_2(matrix_i[178*12+:12]), .o_data(c_plus_d[178][0]), .i_clk(i_clk));
Add0000000001  u_00000000B5_Add0000000001(.i_data_1(matrix_r[179*12+:12]), .i_data_2(matrix_i[179*12+:12]), .o_data(c_plus_d[179][0]), .i_clk(i_clk));
Add0000000001  u_00000000B6_Add0000000001(.i_data_1(matrix_r[180*12+:12]), .i_data_2(matrix_i[180*12+:12]), .o_data(c_plus_d[180][0]), .i_clk(i_clk));
Add0000000001  u_00000000B7_Add0000000001(.i_data_1(matrix_r[181*12+:12]), .i_data_2(matrix_i[181*12+:12]), .o_data(c_plus_d[181][0]), .i_clk(i_clk));
Add0000000001  u_00000000B8_Add0000000001(.i_data_1(matrix_r[182*12+:12]), .i_data_2(matrix_i[182*12+:12]), .o_data(c_plus_d[182][0]), .i_clk(i_clk));
Add0000000001  u_00000000B9_Add0000000001(.i_data_1(matrix_r[183*12+:12]), .i_data_2(matrix_i[183*12+:12]), .o_data(c_plus_d[183][0]), .i_clk(i_clk));
Add0000000001  u_00000000BA_Add0000000001(.i_data_1(matrix_r[184*12+:12]), .i_data_2(matrix_i[184*12+:12]), .o_data(c_plus_d[184][0]), .i_clk(i_clk));
Add0000000001  u_00000000BB_Add0000000001(.i_data_1(matrix_r[185*12+:12]), .i_data_2(matrix_i[185*12+:12]), .o_data(c_plus_d[185][0]), .i_clk(i_clk));
Add0000000001  u_00000000BC_Add0000000001(.i_data_1(matrix_r[186*12+:12]), .i_data_2(matrix_i[186*12+:12]), .o_data(c_plus_d[186][0]), .i_clk(i_clk));
Add0000000001  u_00000000BD_Add0000000001(.i_data_1(matrix_r[187*12+:12]), .i_data_2(matrix_i[187*12+:12]), .o_data(c_plus_d[187][0]), .i_clk(i_clk));
Add0000000001  u_00000000BE_Add0000000001(.i_data_1(matrix_r[188*12+:12]), .i_data_2(matrix_i[188*12+:12]), .o_data(c_plus_d[188][0]), .i_clk(i_clk));
Add0000000001  u_00000000BF_Add0000000001(.i_data_1(matrix_r[189*12+:12]), .i_data_2(matrix_i[189*12+:12]), .o_data(c_plus_d[189][0]), .i_clk(i_clk));
Add0000000001  u_00000000C0_Add0000000001(.i_data_1(matrix_r[190*12+:12]), .i_data_2(matrix_i[190*12+:12]), .o_data(c_plus_d[190][0]), .i_clk(i_clk));
Add0000000001  u_00000000C1_Add0000000001(.i_data_1(matrix_r[191*12+:12]), .i_data_2(matrix_i[191*12+:12]), .o_data(c_plus_d[191][0]), .i_clk(i_clk));
Add0000000001  u_00000000C2_Add0000000001(.i_data_1(matrix_r[192*12+:12]), .i_data_2(matrix_i[192*12+:12]), .o_data(c_plus_d[192][0]), .i_clk(i_clk));
Add0000000001  u_00000000C3_Add0000000001(.i_data_1(matrix_r[193*12+:12]), .i_data_2(matrix_i[193*12+:12]), .o_data(c_plus_d[193][0]), .i_clk(i_clk));
Add0000000001  u_00000000C4_Add0000000001(.i_data_1(matrix_r[194*12+:12]), .i_data_2(matrix_i[194*12+:12]), .o_data(c_plus_d[194][0]), .i_clk(i_clk));
Add0000000001  u_00000000C5_Add0000000001(.i_data_1(matrix_r[195*12+:12]), .i_data_2(matrix_i[195*12+:12]), .o_data(c_plus_d[195][0]), .i_clk(i_clk));
Add0000000001  u_00000000C6_Add0000000001(.i_data_1(matrix_r[196*12+:12]), .i_data_2(matrix_i[196*12+:12]), .o_data(c_plus_d[196][0]), .i_clk(i_clk));
Add0000000001  u_00000000C7_Add0000000001(.i_data_1(matrix_r[197*12+:12]), .i_data_2(matrix_i[197*12+:12]), .o_data(c_plus_d[197][0]), .i_clk(i_clk));
Add0000000001  u_00000000C8_Add0000000001(.i_data_1(matrix_r[198*12+:12]), .i_data_2(matrix_i[198*12+:12]), .o_data(c_plus_d[198][0]), .i_clk(i_clk));
Add0000000001  u_00000000C9_Add0000000001(.i_data_1(matrix_r[199*12+:12]), .i_data_2(matrix_i[199*12+:12]), .o_data(c_plus_d[199][0]), .i_clk(i_clk));
Add0000000001  u_00000000CA_Add0000000001(.i_data_1(matrix_r[200*12+:12]), .i_data_2(matrix_i[200*12+:12]), .o_data(c_plus_d[200][0]), .i_clk(i_clk));
Add0000000001  u_00000000CB_Add0000000001(.i_data_1(matrix_r[201*12+:12]), .i_data_2(matrix_i[201*12+:12]), .o_data(c_plus_d[201][0]), .i_clk(i_clk));
Add0000000001  u_00000000CC_Add0000000001(.i_data_1(matrix_r[202*12+:12]), .i_data_2(matrix_i[202*12+:12]), .o_data(c_plus_d[202][0]), .i_clk(i_clk));
Add0000000001  u_00000000CD_Add0000000001(.i_data_1(matrix_r[203*12+:12]), .i_data_2(matrix_i[203*12+:12]), .o_data(c_plus_d[203][0]), .i_clk(i_clk));
Add0000000001  u_00000000CE_Add0000000001(.i_data_1(matrix_r[204*12+:12]), .i_data_2(matrix_i[204*12+:12]), .o_data(c_plus_d[204][0]), .i_clk(i_clk));
Add0000000001  u_00000000CF_Add0000000001(.i_data_1(matrix_r[205*12+:12]), .i_data_2(matrix_i[205*12+:12]), .o_data(c_plus_d[205][0]), .i_clk(i_clk));
Add0000000001  u_00000000D0_Add0000000001(.i_data_1(matrix_r[206*12+:12]), .i_data_2(matrix_i[206*12+:12]), .o_data(c_plus_d[206][0]), .i_clk(i_clk));
Add0000000001  u_00000000D1_Add0000000001(.i_data_1(matrix_r[207*12+:12]), .i_data_2(matrix_i[207*12+:12]), .o_data(c_plus_d[207][0]), .i_clk(i_clk));
Add0000000001  u_00000000D2_Add0000000001(.i_data_1(matrix_r[208*12+:12]), .i_data_2(matrix_i[208*12+:12]), .o_data(c_plus_d[208][0]), .i_clk(i_clk));
Add0000000001  u_00000000D3_Add0000000001(.i_data_1(matrix_r[209*12+:12]), .i_data_2(matrix_i[209*12+:12]), .o_data(c_plus_d[209][0]), .i_clk(i_clk));
Add0000000001  u_00000000D4_Add0000000001(.i_data_1(matrix_r[210*12+:12]), .i_data_2(matrix_i[210*12+:12]), .o_data(c_plus_d[210][0]), .i_clk(i_clk));
Add0000000001  u_00000000D5_Add0000000001(.i_data_1(matrix_r[211*12+:12]), .i_data_2(matrix_i[211*12+:12]), .o_data(c_plus_d[211][0]), .i_clk(i_clk));
Add0000000001  u_00000000D6_Add0000000001(.i_data_1(matrix_r[212*12+:12]), .i_data_2(matrix_i[212*12+:12]), .o_data(c_plus_d[212][0]), .i_clk(i_clk));
Add0000000001  u_00000000D7_Add0000000001(.i_data_1(matrix_r[213*12+:12]), .i_data_2(matrix_i[213*12+:12]), .o_data(c_plus_d[213][0]), .i_clk(i_clk));
Add0000000001  u_00000000D8_Add0000000001(.i_data_1(matrix_r[214*12+:12]), .i_data_2(matrix_i[214*12+:12]), .o_data(c_plus_d[214][0]), .i_clk(i_clk));
Add0000000001  u_00000000D9_Add0000000001(.i_data_1(matrix_r[215*12+:12]), .i_data_2(matrix_i[215*12+:12]), .o_data(c_plus_d[215][0]), .i_clk(i_clk));
Add0000000001  u_00000000DA_Add0000000001(.i_data_1(matrix_r[216*12+:12]), .i_data_2(matrix_i[216*12+:12]), .o_data(c_plus_d[216][0]), .i_clk(i_clk));
Add0000000001  u_00000000DB_Add0000000001(.i_data_1(matrix_r[217*12+:12]), .i_data_2(matrix_i[217*12+:12]), .o_data(c_plus_d[217][0]), .i_clk(i_clk));
Add0000000001  u_00000000DC_Add0000000001(.i_data_1(matrix_r[218*12+:12]), .i_data_2(matrix_i[218*12+:12]), .o_data(c_plus_d[218][0]), .i_clk(i_clk));
Add0000000001  u_00000000DD_Add0000000001(.i_data_1(matrix_r[219*12+:12]), .i_data_2(matrix_i[219*12+:12]), .o_data(c_plus_d[219][0]), .i_clk(i_clk));
Add0000000001  u_00000000DE_Add0000000001(.i_data_1(matrix_r[220*12+:12]), .i_data_2(matrix_i[220*12+:12]), .o_data(c_plus_d[220][0]), .i_clk(i_clk));
Add0000000001  u_00000000DF_Add0000000001(.i_data_1(matrix_r[221*12+:12]), .i_data_2(matrix_i[221*12+:12]), .o_data(c_plus_d[221][0]), .i_clk(i_clk));
Add0000000001  u_00000000E0_Add0000000001(.i_data_1(matrix_r[222*12+:12]), .i_data_2(matrix_i[222*12+:12]), .o_data(c_plus_d[222][0]), .i_clk(i_clk));
Add0000000001  u_00000000E1_Add0000000001(.i_data_1(matrix_r[223*12+:12]), .i_data_2(matrix_i[223*12+:12]), .o_data(c_plus_d[223][0]), .i_clk(i_clk));
Add0000000001  u_00000000E2_Add0000000001(.i_data_1(matrix_r[224*12+:12]), .i_data_2(matrix_i[224*12+:12]), .o_data(c_plus_d[224][0]), .i_clk(i_clk));
Add0000000001  u_00000000E3_Add0000000001(.i_data_1(matrix_r[225*12+:12]), .i_data_2(matrix_i[225*12+:12]), .o_data(c_plus_d[225][0]), .i_clk(i_clk));
Add0000000001  u_00000000E4_Add0000000001(.i_data_1(matrix_r[226*12+:12]), .i_data_2(matrix_i[226*12+:12]), .o_data(c_plus_d[226][0]), .i_clk(i_clk));
Add0000000001  u_00000000E5_Add0000000001(.i_data_1(matrix_r[227*12+:12]), .i_data_2(matrix_i[227*12+:12]), .o_data(c_plus_d[227][0]), .i_clk(i_clk));
Add0000000001  u_00000000E6_Add0000000001(.i_data_1(matrix_r[228*12+:12]), .i_data_2(matrix_i[228*12+:12]), .o_data(c_plus_d[228][0]), .i_clk(i_clk));
Add0000000001  u_00000000E7_Add0000000001(.i_data_1(matrix_r[229*12+:12]), .i_data_2(matrix_i[229*12+:12]), .o_data(c_plus_d[229][0]), .i_clk(i_clk));
Add0000000001  u_00000000E8_Add0000000001(.i_data_1(matrix_r[230*12+:12]), .i_data_2(matrix_i[230*12+:12]), .o_data(c_plus_d[230][0]), .i_clk(i_clk));
Add0000000001  u_00000000E9_Add0000000001(.i_data_1(matrix_r[231*12+:12]), .i_data_2(matrix_i[231*12+:12]), .o_data(c_plus_d[231][0]), .i_clk(i_clk));
Add0000000001  u_00000000EA_Add0000000001(.i_data_1(matrix_r[232*12+:12]), .i_data_2(matrix_i[232*12+:12]), .o_data(c_plus_d[232][0]), .i_clk(i_clk));
Add0000000001  u_00000000EB_Add0000000001(.i_data_1(matrix_r[233*12+:12]), .i_data_2(matrix_i[233*12+:12]), .o_data(c_plus_d[233][0]), .i_clk(i_clk));
Add0000000001  u_00000000EC_Add0000000001(.i_data_1(matrix_r[234*12+:12]), .i_data_2(matrix_i[234*12+:12]), .o_data(c_plus_d[234][0]), .i_clk(i_clk));
Add0000000001  u_00000000ED_Add0000000001(.i_data_1(matrix_r[235*12+:12]), .i_data_2(matrix_i[235*12+:12]), .o_data(c_plus_d[235][0]), .i_clk(i_clk));
Add0000000001  u_00000000EE_Add0000000001(.i_data_1(matrix_r[236*12+:12]), .i_data_2(matrix_i[236*12+:12]), .o_data(c_plus_d[236][0]), .i_clk(i_clk));
Add0000000001  u_00000000EF_Add0000000001(.i_data_1(matrix_r[237*12+:12]), .i_data_2(matrix_i[237*12+:12]), .o_data(c_plus_d[237][0]), .i_clk(i_clk));
Add0000000001  u_00000000F0_Add0000000001(.i_data_1(matrix_r[238*12+:12]), .i_data_2(matrix_i[238*12+:12]), .o_data(c_plus_d[238][0]), .i_clk(i_clk));
Add0000000001  u_00000000F1_Add0000000001(.i_data_1(matrix_r[239*12+:12]), .i_data_2(matrix_i[239*12+:12]), .o_data(c_plus_d[239][0]), .i_clk(i_clk));
Add0000000001  u_00000000F2_Add0000000001(.i_data_1(matrix_r[240*12+:12]), .i_data_2(matrix_i[240*12+:12]), .o_data(c_plus_d[240][0]), .i_clk(i_clk));
Add0000000001  u_00000000F3_Add0000000001(.i_data_1(matrix_r[241*12+:12]), .i_data_2(matrix_i[241*12+:12]), .o_data(c_plus_d[241][0]), .i_clk(i_clk));
Add0000000001  u_00000000F4_Add0000000001(.i_data_1(matrix_r[242*12+:12]), .i_data_2(matrix_i[242*12+:12]), .o_data(c_plus_d[242][0]), .i_clk(i_clk));
Add0000000001  u_00000000F5_Add0000000001(.i_data_1(matrix_r[243*12+:12]), .i_data_2(matrix_i[243*12+:12]), .o_data(c_plus_d[243][0]), .i_clk(i_clk));
Add0000000001  u_00000000F6_Add0000000001(.i_data_1(matrix_r[244*12+:12]), .i_data_2(matrix_i[244*12+:12]), .o_data(c_plus_d[244][0]), .i_clk(i_clk));
Add0000000001  u_00000000F7_Add0000000001(.i_data_1(matrix_r[245*12+:12]), .i_data_2(matrix_i[245*12+:12]), .o_data(c_plus_d[245][0]), .i_clk(i_clk));
Add0000000001  u_00000000F8_Add0000000001(.i_data_1(matrix_r[246*12+:12]), .i_data_2(matrix_i[246*12+:12]), .o_data(c_plus_d[246][0]), .i_clk(i_clk));
Add0000000001  u_00000000F9_Add0000000001(.i_data_1(matrix_r[247*12+:12]), .i_data_2(matrix_i[247*12+:12]), .o_data(c_plus_d[247][0]), .i_clk(i_clk));
Add0000000001  u_00000000FA_Add0000000001(.i_data_1(matrix_r[248*12+:12]), .i_data_2(matrix_i[248*12+:12]), .o_data(c_plus_d[248][0]), .i_clk(i_clk));
Add0000000001  u_00000000FB_Add0000000001(.i_data_1(matrix_r[249*12+:12]), .i_data_2(matrix_i[249*12+:12]), .o_data(c_plus_d[249][0]), .i_clk(i_clk));
Add0000000001  u_00000000FC_Add0000000001(.i_data_1(matrix_r[250*12+:12]), .i_data_2(matrix_i[250*12+:12]), .o_data(c_plus_d[250][0]), .i_clk(i_clk));
Add0000000001  u_00000000FD_Add0000000001(.i_data_1(matrix_r[251*12+:12]), .i_data_2(matrix_i[251*12+:12]), .o_data(c_plus_d[251][0]), .i_clk(i_clk));
Add0000000001  u_00000000FE_Add0000000001(.i_data_1(matrix_r[252*12+:12]), .i_data_2(matrix_i[252*12+:12]), .o_data(c_plus_d[252][0]), .i_clk(i_clk));
Add0000000001  u_00000000FF_Add0000000001(.i_data_1(matrix_r[253*12+:12]), .i_data_2(matrix_i[253*12+:12]), .o_data(c_plus_d[253][0]), .i_clk(i_clk));
Add0000000001  u_0000000100_Add0000000001(.i_data_1(matrix_r[254*12+:12]), .i_data_2(matrix_i[254*12+:12]), .o_data(c_plus_d[254][0]), .i_clk(i_clk));
Add0000000001  u_0000000101_Add0000000001(.i_data_1(matrix_r[255*12+:12]), .i_data_2(matrix_i[255*12+:12]), .o_data(c_plus_d[255][0]), .i_clk(i_clk));
Add0000000001  u_0000000102_Add0000000001(.i_data_1(vector_r[1*12+:12]), .i_data_2(vector_i[1*12+:12]), .o_data(a_plus_b[1]), .i_clk(i_clk));
Sub0000000001  u_0000000002_Sub0000000001(.i_data_1(vector_i[1*12+:12]), .i_data_2(vector_r[1*12+:12]), .o_data(b_minus_a[1]), .i_clk(i_clk));
Add0000000001  u_0000000103_Add0000000001(.i_data_1(matrix_r[256*12+:12]), .i_data_2(matrix_i[256*12+:12]), .o_data(c_plus_d[0][1]), .i_clk(i_clk));
Add0000000001  u_0000000104_Add0000000001(.i_data_1(matrix_r[257*12+:12]), .i_data_2(matrix_i[257*12+:12]), .o_data(c_plus_d[1][1]), .i_clk(i_clk));
Add0000000001  u_0000000105_Add0000000001(.i_data_1(matrix_r[258*12+:12]), .i_data_2(matrix_i[258*12+:12]), .o_data(c_plus_d[2][1]), .i_clk(i_clk));
Add0000000001  u_0000000106_Add0000000001(.i_data_1(matrix_r[259*12+:12]), .i_data_2(matrix_i[259*12+:12]), .o_data(c_plus_d[3][1]), .i_clk(i_clk));
Add0000000001  u_0000000107_Add0000000001(.i_data_1(matrix_r[260*12+:12]), .i_data_2(matrix_i[260*12+:12]), .o_data(c_plus_d[4][1]), .i_clk(i_clk));
Add0000000001  u_0000000108_Add0000000001(.i_data_1(matrix_r[261*12+:12]), .i_data_2(matrix_i[261*12+:12]), .o_data(c_plus_d[5][1]), .i_clk(i_clk));
Add0000000001  u_0000000109_Add0000000001(.i_data_1(matrix_r[262*12+:12]), .i_data_2(matrix_i[262*12+:12]), .o_data(c_plus_d[6][1]), .i_clk(i_clk));
Add0000000001  u_000000010A_Add0000000001(.i_data_1(matrix_r[263*12+:12]), .i_data_2(matrix_i[263*12+:12]), .o_data(c_plus_d[7][1]), .i_clk(i_clk));
Add0000000001  u_000000010B_Add0000000001(.i_data_1(matrix_r[264*12+:12]), .i_data_2(matrix_i[264*12+:12]), .o_data(c_plus_d[8][1]), .i_clk(i_clk));
Add0000000001  u_000000010C_Add0000000001(.i_data_1(matrix_r[265*12+:12]), .i_data_2(matrix_i[265*12+:12]), .o_data(c_plus_d[9][1]), .i_clk(i_clk));
Add0000000001  u_000000010D_Add0000000001(.i_data_1(matrix_r[266*12+:12]), .i_data_2(matrix_i[266*12+:12]), .o_data(c_plus_d[10][1]), .i_clk(i_clk));
Add0000000001  u_000000010E_Add0000000001(.i_data_1(matrix_r[267*12+:12]), .i_data_2(matrix_i[267*12+:12]), .o_data(c_plus_d[11][1]), .i_clk(i_clk));
Add0000000001  u_000000010F_Add0000000001(.i_data_1(matrix_r[268*12+:12]), .i_data_2(matrix_i[268*12+:12]), .o_data(c_plus_d[12][1]), .i_clk(i_clk));
Add0000000001  u_0000000110_Add0000000001(.i_data_1(matrix_r[269*12+:12]), .i_data_2(matrix_i[269*12+:12]), .o_data(c_plus_d[13][1]), .i_clk(i_clk));
Add0000000001  u_0000000111_Add0000000001(.i_data_1(matrix_r[270*12+:12]), .i_data_2(matrix_i[270*12+:12]), .o_data(c_plus_d[14][1]), .i_clk(i_clk));
Add0000000001  u_0000000112_Add0000000001(.i_data_1(matrix_r[271*12+:12]), .i_data_2(matrix_i[271*12+:12]), .o_data(c_plus_d[15][1]), .i_clk(i_clk));
Add0000000001  u_0000000113_Add0000000001(.i_data_1(matrix_r[272*12+:12]), .i_data_2(matrix_i[272*12+:12]), .o_data(c_plus_d[16][1]), .i_clk(i_clk));
Add0000000001  u_0000000114_Add0000000001(.i_data_1(matrix_r[273*12+:12]), .i_data_2(matrix_i[273*12+:12]), .o_data(c_plus_d[17][1]), .i_clk(i_clk));
Add0000000001  u_0000000115_Add0000000001(.i_data_1(matrix_r[274*12+:12]), .i_data_2(matrix_i[274*12+:12]), .o_data(c_plus_d[18][1]), .i_clk(i_clk));
Add0000000001  u_0000000116_Add0000000001(.i_data_1(matrix_r[275*12+:12]), .i_data_2(matrix_i[275*12+:12]), .o_data(c_plus_d[19][1]), .i_clk(i_clk));
Add0000000001  u_0000000117_Add0000000001(.i_data_1(matrix_r[276*12+:12]), .i_data_2(matrix_i[276*12+:12]), .o_data(c_plus_d[20][1]), .i_clk(i_clk));
Add0000000001  u_0000000118_Add0000000001(.i_data_1(matrix_r[277*12+:12]), .i_data_2(matrix_i[277*12+:12]), .o_data(c_plus_d[21][1]), .i_clk(i_clk));
Add0000000001  u_0000000119_Add0000000001(.i_data_1(matrix_r[278*12+:12]), .i_data_2(matrix_i[278*12+:12]), .o_data(c_plus_d[22][1]), .i_clk(i_clk));
Add0000000001  u_000000011A_Add0000000001(.i_data_1(matrix_r[279*12+:12]), .i_data_2(matrix_i[279*12+:12]), .o_data(c_plus_d[23][1]), .i_clk(i_clk));
Add0000000001  u_000000011B_Add0000000001(.i_data_1(matrix_r[280*12+:12]), .i_data_2(matrix_i[280*12+:12]), .o_data(c_plus_d[24][1]), .i_clk(i_clk));
Add0000000001  u_000000011C_Add0000000001(.i_data_1(matrix_r[281*12+:12]), .i_data_2(matrix_i[281*12+:12]), .o_data(c_plus_d[25][1]), .i_clk(i_clk));
Add0000000001  u_000000011D_Add0000000001(.i_data_1(matrix_r[282*12+:12]), .i_data_2(matrix_i[282*12+:12]), .o_data(c_plus_d[26][1]), .i_clk(i_clk));
Add0000000001  u_000000011E_Add0000000001(.i_data_1(matrix_r[283*12+:12]), .i_data_2(matrix_i[283*12+:12]), .o_data(c_plus_d[27][1]), .i_clk(i_clk));
Add0000000001  u_000000011F_Add0000000001(.i_data_1(matrix_r[284*12+:12]), .i_data_2(matrix_i[284*12+:12]), .o_data(c_plus_d[28][1]), .i_clk(i_clk));
Add0000000001  u_0000000120_Add0000000001(.i_data_1(matrix_r[285*12+:12]), .i_data_2(matrix_i[285*12+:12]), .o_data(c_plus_d[29][1]), .i_clk(i_clk));
Add0000000001  u_0000000121_Add0000000001(.i_data_1(matrix_r[286*12+:12]), .i_data_2(matrix_i[286*12+:12]), .o_data(c_plus_d[30][1]), .i_clk(i_clk));
Add0000000001  u_0000000122_Add0000000001(.i_data_1(matrix_r[287*12+:12]), .i_data_2(matrix_i[287*12+:12]), .o_data(c_plus_d[31][1]), .i_clk(i_clk));
Add0000000001  u_0000000123_Add0000000001(.i_data_1(matrix_r[288*12+:12]), .i_data_2(matrix_i[288*12+:12]), .o_data(c_plus_d[32][1]), .i_clk(i_clk));
Add0000000001  u_0000000124_Add0000000001(.i_data_1(matrix_r[289*12+:12]), .i_data_2(matrix_i[289*12+:12]), .o_data(c_plus_d[33][1]), .i_clk(i_clk));
Add0000000001  u_0000000125_Add0000000001(.i_data_1(matrix_r[290*12+:12]), .i_data_2(matrix_i[290*12+:12]), .o_data(c_plus_d[34][1]), .i_clk(i_clk));
Add0000000001  u_0000000126_Add0000000001(.i_data_1(matrix_r[291*12+:12]), .i_data_2(matrix_i[291*12+:12]), .o_data(c_plus_d[35][1]), .i_clk(i_clk));
Add0000000001  u_0000000127_Add0000000001(.i_data_1(matrix_r[292*12+:12]), .i_data_2(matrix_i[292*12+:12]), .o_data(c_plus_d[36][1]), .i_clk(i_clk));
Add0000000001  u_0000000128_Add0000000001(.i_data_1(matrix_r[293*12+:12]), .i_data_2(matrix_i[293*12+:12]), .o_data(c_plus_d[37][1]), .i_clk(i_clk));
Add0000000001  u_0000000129_Add0000000001(.i_data_1(matrix_r[294*12+:12]), .i_data_2(matrix_i[294*12+:12]), .o_data(c_plus_d[38][1]), .i_clk(i_clk));
Add0000000001  u_000000012A_Add0000000001(.i_data_1(matrix_r[295*12+:12]), .i_data_2(matrix_i[295*12+:12]), .o_data(c_plus_d[39][1]), .i_clk(i_clk));
Add0000000001  u_000000012B_Add0000000001(.i_data_1(matrix_r[296*12+:12]), .i_data_2(matrix_i[296*12+:12]), .o_data(c_plus_d[40][1]), .i_clk(i_clk));
Add0000000001  u_000000012C_Add0000000001(.i_data_1(matrix_r[297*12+:12]), .i_data_2(matrix_i[297*12+:12]), .o_data(c_plus_d[41][1]), .i_clk(i_clk));
Add0000000001  u_000000012D_Add0000000001(.i_data_1(matrix_r[298*12+:12]), .i_data_2(matrix_i[298*12+:12]), .o_data(c_plus_d[42][1]), .i_clk(i_clk));
Add0000000001  u_000000012E_Add0000000001(.i_data_1(matrix_r[299*12+:12]), .i_data_2(matrix_i[299*12+:12]), .o_data(c_plus_d[43][1]), .i_clk(i_clk));
Add0000000001  u_000000012F_Add0000000001(.i_data_1(matrix_r[300*12+:12]), .i_data_2(matrix_i[300*12+:12]), .o_data(c_plus_d[44][1]), .i_clk(i_clk));
Add0000000001  u_0000000130_Add0000000001(.i_data_1(matrix_r[301*12+:12]), .i_data_2(matrix_i[301*12+:12]), .o_data(c_plus_d[45][1]), .i_clk(i_clk));
Add0000000001  u_0000000131_Add0000000001(.i_data_1(matrix_r[302*12+:12]), .i_data_2(matrix_i[302*12+:12]), .o_data(c_plus_d[46][1]), .i_clk(i_clk));
Add0000000001  u_0000000132_Add0000000001(.i_data_1(matrix_r[303*12+:12]), .i_data_2(matrix_i[303*12+:12]), .o_data(c_plus_d[47][1]), .i_clk(i_clk));
Add0000000001  u_0000000133_Add0000000001(.i_data_1(matrix_r[304*12+:12]), .i_data_2(matrix_i[304*12+:12]), .o_data(c_plus_d[48][1]), .i_clk(i_clk));
Add0000000001  u_0000000134_Add0000000001(.i_data_1(matrix_r[305*12+:12]), .i_data_2(matrix_i[305*12+:12]), .o_data(c_plus_d[49][1]), .i_clk(i_clk));
Add0000000001  u_0000000135_Add0000000001(.i_data_1(matrix_r[306*12+:12]), .i_data_2(matrix_i[306*12+:12]), .o_data(c_plus_d[50][1]), .i_clk(i_clk));
Add0000000001  u_0000000136_Add0000000001(.i_data_1(matrix_r[307*12+:12]), .i_data_2(matrix_i[307*12+:12]), .o_data(c_plus_d[51][1]), .i_clk(i_clk));
Add0000000001  u_0000000137_Add0000000001(.i_data_1(matrix_r[308*12+:12]), .i_data_2(matrix_i[308*12+:12]), .o_data(c_plus_d[52][1]), .i_clk(i_clk));
Add0000000001  u_0000000138_Add0000000001(.i_data_1(matrix_r[309*12+:12]), .i_data_2(matrix_i[309*12+:12]), .o_data(c_plus_d[53][1]), .i_clk(i_clk));
Add0000000001  u_0000000139_Add0000000001(.i_data_1(matrix_r[310*12+:12]), .i_data_2(matrix_i[310*12+:12]), .o_data(c_plus_d[54][1]), .i_clk(i_clk));
Add0000000001  u_000000013A_Add0000000001(.i_data_1(matrix_r[311*12+:12]), .i_data_2(matrix_i[311*12+:12]), .o_data(c_plus_d[55][1]), .i_clk(i_clk));
Add0000000001  u_000000013B_Add0000000001(.i_data_1(matrix_r[312*12+:12]), .i_data_2(matrix_i[312*12+:12]), .o_data(c_plus_d[56][1]), .i_clk(i_clk));
Add0000000001  u_000000013C_Add0000000001(.i_data_1(matrix_r[313*12+:12]), .i_data_2(matrix_i[313*12+:12]), .o_data(c_plus_d[57][1]), .i_clk(i_clk));
Add0000000001  u_000000013D_Add0000000001(.i_data_1(matrix_r[314*12+:12]), .i_data_2(matrix_i[314*12+:12]), .o_data(c_plus_d[58][1]), .i_clk(i_clk));
Add0000000001  u_000000013E_Add0000000001(.i_data_1(matrix_r[315*12+:12]), .i_data_2(matrix_i[315*12+:12]), .o_data(c_plus_d[59][1]), .i_clk(i_clk));
Add0000000001  u_000000013F_Add0000000001(.i_data_1(matrix_r[316*12+:12]), .i_data_2(matrix_i[316*12+:12]), .o_data(c_plus_d[60][1]), .i_clk(i_clk));
Add0000000001  u_0000000140_Add0000000001(.i_data_1(matrix_r[317*12+:12]), .i_data_2(matrix_i[317*12+:12]), .o_data(c_plus_d[61][1]), .i_clk(i_clk));
Add0000000001  u_0000000141_Add0000000001(.i_data_1(matrix_r[318*12+:12]), .i_data_2(matrix_i[318*12+:12]), .o_data(c_plus_d[62][1]), .i_clk(i_clk));
Add0000000001  u_0000000142_Add0000000001(.i_data_1(matrix_r[319*12+:12]), .i_data_2(matrix_i[319*12+:12]), .o_data(c_plus_d[63][1]), .i_clk(i_clk));
Add0000000001  u_0000000143_Add0000000001(.i_data_1(matrix_r[320*12+:12]), .i_data_2(matrix_i[320*12+:12]), .o_data(c_plus_d[64][1]), .i_clk(i_clk));
Add0000000001  u_0000000144_Add0000000001(.i_data_1(matrix_r[321*12+:12]), .i_data_2(matrix_i[321*12+:12]), .o_data(c_plus_d[65][1]), .i_clk(i_clk));
Add0000000001  u_0000000145_Add0000000001(.i_data_1(matrix_r[322*12+:12]), .i_data_2(matrix_i[322*12+:12]), .o_data(c_plus_d[66][1]), .i_clk(i_clk));
Add0000000001  u_0000000146_Add0000000001(.i_data_1(matrix_r[323*12+:12]), .i_data_2(matrix_i[323*12+:12]), .o_data(c_plus_d[67][1]), .i_clk(i_clk));
Add0000000001  u_0000000147_Add0000000001(.i_data_1(matrix_r[324*12+:12]), .i_data_2(matrix_i[324*12+:12]), .o_data(c_plus_d[68][1]), .i_clk(i_clk));
Add0000000001  u_0000000148_Add0000000001(.i_data_1(matrix_r[325*12+:12]), .i_data_2(matrix_i[325*12+:12]), .o_data(c_plus_d[69][1]), .i_clk(i_clk));
Add0000000001  u_0000000149_Add0000000001(.i_data_1(matrix_r[326*12+:12]), .i_data_2(matrix_i[326*12+:12]), .o_data(c_plus_d[70][1]), .i_clk(i_clk));
Add0000000001  u_000000014A_Add0000000001(.i_data_1(matrix_r[327*12+:12]), .i_data_2(matrix_i[327*12+:12]), .o_data(c_plus_d[71][1]), .i_clk(i_clk));
Add0000000001  u_000000014B_Add0000000001(.i_data_1(matrix_r[328*12+:12]), .i_data_2(matrix_i[328*12+:12]), .o_data(c_plus_d[72][1]), .i_clk(i_clk));
Add0000000001  u_000000014C_Add0000000001(.i_data_1(matrix_r[329*12+:12]), .i_data_2(matrix_i[329*12+:12]), .o_data(c_plus_d[73][1]), .i_clk(i_clk));
Add0000000001  u_000000014D_Add0000000001(.i_data_1(matrix_r[330*12+:12]), .i_data_2(matrix_i[330*12+:12]), .o_data(c_plus_d[74][1]), .i_clk(i_clk));
Add0000000001  u_000000014E_Add0000000001(.i_data_1(matrix_r[331*12+:12]), .i_data_2(matrix_i[331*12+:12]), .o_data(c_plus_d[75][1]), .i_clk(i_clk));
Add0000000001  u_000000014F_Add0000000001(.i_data_1(matrix_r[332*12+:12]), .i_data_2(matrix_i[332*12+:12]), .o_data(c_plus_d[76][1]), .i_clk(i_clk));
Add0000000001  u_0000000150_Add0000000001(.i_data_1(matrix_r[333*12+:12]), .i_data_2(matrix_i[333*12+:12]), .o_data(c_plus_d[77][1]), .i_clk(i_clk));
Add0000000001  u_0000000151_Add0000000001(.i_data_1(matrix_r[334*12+:12]), .i_data_2(matrix_i[334*12+:12]), .o_data(c_plus_d[78][1]), .i_clk(i_clk));
Add0000000001  u_0000000152_Add0000000001(.i_data_1(matrix_r[335*12+:12]), .i_data_2(matrix_i[335*12+:12]), .o_data(c_plus_d[79][1]), .i_clk(i_clk));
Add0000000001  u_0000000153_Add0000000001(.i_data_1(matrix_r[336*12+:12]), .i_data_2(matrix_i[336*12+:12]), .o_data(c_plus_d[80][1]), .i_clk(i_clk));
Add0000000001  u_0000000154_Add0000000001(.i_data_1(matrix_r[337*12+:12]), .i_data_2(matrix_i[337*12+:12]), .o_data(c_plus_d[81][1]), .i_clk(i_clk));
Add0000000001  u_0000000155_Add0000000001(.i_data_1(matrix_r[338*12+:12]), .i_data_2(matrix_i[338*12+:12]), .o_data(c_plus_d[82][1]), .i_clk(i_clk));
Add0000000001  u_0000000156_Add0000000001(.i_data_1(matrix_r[339*12+:12]), .i_data_2(matrix_i[339*12+:12]), .o_data(c_plus_d[83][1]), .i_clk(i_clk));
Add0000000001  u_0000000157_Add0000000001(.i_data_1(matrix_r[340*12+:12]), .i_data_2(matrix_i[340*12+:12]), .o_data(c_plus_d[84][1]), .i_clk(i_clk));
Add0000000001  u_0000000158_Add0000000001(.i_data_1(matrix_r[341*12+:12]), .i_data_2(matrix_i[341*12+:12]), .o_data(c_plus_d[85][1]), .i_clk(i_clk));
Add0000000001  u_0000000159_Add0000000001(.i_data_1(matrix_r[342*12+:12]), .i_data_2(matrix_i[342*12+:12]), .o_data(c_plus_d[86][1]), .i_clk(i_clk));
Add0000000001  u_000000015A_Add0000000001(.i_data_1(matrix_r[343*12+:12]), .i_data_2(matrix_i[343*12+:12]), .o_data(c_plus_d[87][1]), .i_clk(i_clk));
Add0000000001  u_000000015B_Add0000000001(.i_data_1(matrix_r[344*12+:12]), .i_data_2(matrix_i[344*12+:12]), .o_data(c_plus_d[88][1]), .i_clk(i_clk));
Add0000000001  u_000000015C_Add0000000001(.i_data_1(matrix_r[345*12+:12]), .i_data_2(matrix_i[345*12+:12]), .o_data(c_plus_d[89][1]), .i_clk(i_clk));
Add0000000001  u_000000015D_Add0000000001(.i_data_1(matrix_r[346*12+:12]), .i_data_2(matrix_i[346*12+:12]), .o_data(c_plus_d[90][1]), .i_clk(i_clk));
Add0000000001  u_000000015E_Add0000000001(.i_data_1(matrix_r[347*12+:12]), .i_data_2(matrix_i[347*12+:12]), .o_data(c_plus_d[91][1]), .i_clk(i_clk));
Add0000000001  u_000000015F_Add0000000001(.i_data_1(matrix_r[348*12+:12]), .i_data_2(matrix_i[348*12+:12]), .o_data(c_plus_d[92][1]), .i_clk(i_clk));
Add0000000001  u_0000000160_Add0000000001(.i_data_1(matrix_r[349*12+:12]), .i_data_2(matrix_i[349*12+:12]), .o_data(c_plus_d[93][1]), .i_clk(i_clk));
Add0000000001  u_0000000161_Add0000000001(.i_data_1(matrix_r[350*12+:12]), .i_data_2(matrix_i[350*12+:12]), .o_data(c_plus_d[94][1]), .i_clk(i_clk));
Add0000000001  u_0000000162_Add0000000001(.i_data_1(matrix_r[351*12+:12]), .i_data_2(matrix_i[351*12+:12]), .o_data(c_plus_d[95][1]), .i_clk(i_clk));
Add0000000001  u_0000000163_Add0000000001(.i_data_1(matrix_r[352*12+:12]), .i_data_2(matrix_i[352*12+:12]), .o_data(c_plus_d[96][1]), .i_clk(i_clk));
Add0000000001  u_0000000164_Add0000000001(.i_data_1(matrix_r[353*12+:12]), .i_data_2(matrix_i[353*12+:12]), .o_data(c_plus_d[97][1]), .i_clk(i_clk));
Add0000000001  u_0000000165_Add0000000001(.i_data_1(matrix_r[354*12+:12]), .i_data_2(matrix_i[354*12+:12]), .o_data(c_plus_d[98][1]), .i_clk(i_clk));
Add0000000001  u_0000000166_Add0000000001(.i_data_1(matrix_r[355*12+:12]), .i_data_2(matrix_i[355*12+:12]), .o_data(c_plus_d[99][1]), .i_clk(i_clk));
Add0000000001  u_0000000167_Add0000000001(.i_data_1(matrix_r[356*12+:12]), .i_data_2(matrix_i[356*12+:12]), .o_data(c_plus_d[100][1]), .i_clk(i_clk));
Add0000000001  u_0000000168_Add0000000001(.i_data_1(matrix_r[357*12+:12]), .i_data_2(matrix_i[357*12+:12]), .o_data(c_plus_d[101][1]), .i_clk(i_clk));
Add0000000001  u_0000000169_Add0000000001(.i_data_1(matrix_r[358*12+:12]), .i_data_2(matrix_i[358*12+:12]), .o_data(c_plus_d[102][1]), .i_clk(i_clk));
Add0000000001  u_000000016A_Add0000000001(.i_data_1(matrix_r[359*12+:12]), .i_data_2(matrix_i[359*12+:12]), .o_data(c_plus_d[103][1]), .i_clk(i_clk));
Add0000000001  u_000000016B_Add0000000001(.i_data_1(matrix_r[360*12+:12]), .i_data_2(matrix_i[360*12+:12]), .o_data(c_plus_d[104][1]), .i_clk(i_clk));
Add0000000001  u_000000016C_Add0000000001(.i_data_1(matrix_r[361*12+:12]), .i_data_2(matrix_i[361*12+:12]), .o_data(c_plus_d[105][1]), .i_clk(i_clk));
Add0000000001  u_000000016D_Add0000000001(.i_data_1(matrix_r[362*12+:12]), .i_data_2(matrix_i[362*12+:12]), .o_data(c_plus_d[106][1]), .i_clk(i_clk));
Add0000000001  u_000000016E_Add0000000001(.i_data_1(matrix_r[363*12+:12]), .i_data_2(matrix_i[363*12+:12]), .o_data(c_plus_d[107][1]), .i_clk(i_clk));
Add0000000001  u_000000016F_Add0000000001(.i_data_1(matrix_r[364*12+:12]), .i_data_2(matrix_i[364*12+:12]), .o_data(c_plus_d[108][1]), .i_clk(i_clk));
Add0000000001  u_0000000170_Add0000000001(.i_data_1(matrix_r[365*12+:12]), .i_data_2(matrix_i[365*12+:12]), .o_data(c_plus_d[109][1]), .i_clk(i_clk));
Add0000000001  u_0000000171_Add0000000001(.i_data_1(matrix_r[366*12+:12]), .i_data_2(matrix_i[366*12+:12]), .o_data(c_plus_d[110][1]), .i_clk(i_clk));
Add0000000001  u_0000000172_Add0000000001(.i_data_1(matrix_r[367*12+:12]), .i_data_2(matrix_i[367*12+:12]), .o_data(c_plus_d[111][1]), .i_clk(i_clk));
Add0000000001  u_0000000173_Add0000000001(.i_data_1(matrix_r[368*12+:12]), .i_data_2(matrix_i[368*12+:12]), .o_data(c_plus_d[112][1]), .i_clk(i_clk));
Add0000000001  u_0000000174_Add0000000001(.i_data_1(matrix_r[369*12+:12]), .i_data_2(matrix_i[369*12+:12]), .o_data(c_plus_d[113][1]), .i_clk(i_clk));
Add0000000001  u_0000000175_Add0000000001(.i_data_1(matrix_r[370*12+:12]), .i_data_2(matrix_i[370*12+:12]), .o_data(c_plus_d[114][1]), .i_clk(i_clk));
Add0000000001  u_0000000176_Add0000000001(.i_data_1(matrix_r[371*12+:12]), .i_data_2(matrix_i[371*12+:12]), .o_data(c_plus_d[115][1]), .i_clk(i_clk));
Add0000000001  u_0000000177_Add0000000001(.i_data_1(matrix_r[372*12+:12]), .i_data_2(matrix_i[372*12+:12]), .o_data(c_plus_d[116][1]), .i_clk(i_clk));
Add0000000001  u_0000000178_Add0000000001(.i_data_1(matrix_r[373*12+:12]), .i_data_2(matrix_i[373*12+:12]), .o_data(c_plus_d[117][1]), .i_clk(i_clk));
Add0000000001  u_0000000179_Add0000000001(.i_data_1(matrix_r[374*12+:12]), .i_data_2(matrix_i[374*12+:12]), .o_data(c_plus_d[118][1]), .i_clk(i_clk));
Add0000000001  u_000000017A_Add0000000001(.i_data_1(matrix_r[375*12+:12]), .i_data_2(matrix_i[375*12+:12]), .o_data(c_plus_d[119][1]), .i_clk(i_clk));
Add0000000001  u_000000017B_Add0000000001(.i_data_1(matrix_r[376*12+:12]), .i_data_2(matrix_i[376*12+:12]), .o_data(c_plus_d[120][1]), .i_clk(i_clk));
Add0000000001  u_000000017C_Add0000000001(.i_data_1(matrix_r[377*12+:12]), .i_data_2(matrix_i[377*12+:12]), .o_data(c_plus_d[121][1]), .i_clk(i_clk));
Add0000000001  u_000000017D_Add0000000001(.i_data_1(matrix_r[378*12+:12]), .i_data_2(matrix_i[378*12+:12]), .o_data(c_plus_d[122][1]), .i_clk(i_clk));
Add0000000001  u_000000017E_Add0000000001(.i_data_1(matrix_r[379*12+:12]), .i_data_2(matrix_i[379*12+:12]), .o_data(c_plus_d[123][1]), .i_clk(i_clk));
Add0000000001  u_000000017F_Add0000000001(.i_data_1(matrix_r[380*12+:12]), .i_data_2(matrix_i[380*12+:12]), .o_data(c_plus_d[124][1]), .i_clk(i_clk));
Add0000000001  u_0000000180_Add0000000001(.i_data_1(matrix_r[381*12+:12]), .i_data_2(matrix_i[381*12+:12]), .o_data(c_plus_d[125][1]), .i_clk(i_clk));
Add0000000001  u_0000000181_Add0000000001(.i_data_1(matrix_r[382*12+:12]), .i_data_2(matrix_i[382*12+:12]), .o_data(c_plus_d[126][1]), .i_clk(i_clk));
Add0000000001  u_0000000182_Add0000000001(.i_data_1(matrix_r[383*12+:12]), .i_data_2(matrix_i[383*12+:12]), .o_data(c_plus_d[127][1]), .i_clk(i_clk));
Add0000000001  u_0000000183_Add0000000001(.i_data_1(matrix_r[384*12+:12]), .i_data_2(matrix_i[384*12+:12]), .o_data(c_plus_d[128][1]), .i_clk(i_clk));
Add0000000001  u_0000000184_Add0000000001(.i_data_1(matrix_r[385*12+:12]), .i_data_2(matrix_i[385*12+:12]), .o_data(c_plus_d[129][1]), .i_clk(i_clk));
Add0000000001  u_0000000185_Add0000000001(.i_data_1(matrix_r[386*12+:12]), .i_data_2(matrix_i[386*12+:12]), .o_data(c_plus_d[130][1]), .i_clk(i_clk));
Add0000000001  u_0000000186_Add0000000001(.i_data_1(matrix_r[387*12+:12]), .i_data_2(matrix_i[387*12+:12]), .o_data(c_plus_d[131][1]), .i_clk(i_clk));
Add0000000001  u_0000000187_Add0000000001(.i_data_1(matrix_r[388*12+:12]), .i_data_2(matrix_i[388*12+:12]), .o_data(c_plus_d[132][1]), .i_clk(i_clk));
Add0000000001  u_0000000188_Add0000000001(.i_data_1(matrix_r[389*12+:12]), .i_data_2(matrix_i[389*12+:12]), .o_data(c_plus_d[133][1]), .i_clk(i_clk));
Add0000000001  u_0000000189_Add0000000001(.i_data_1(matrix_r[390*12+:12]), .i_data_2(matrix_i[390*12+:12]), .o_data(c_plus_d[134][1]), .i_clk(i_clk));
Add0000000001  u_000000018A_Add0000000001(.i_data_1(matrix_r[391*12+:12]), .i_data_2(matrix_i[391*12+:12]), .o_data(c_plus_d[135][1]), .i_clk(i_clk));
Add0000000001  u_000000018B_Add0000000001(.i_data_1(matrix_r[392*12+:12]), .i_data_2(matrix_i[392*12+:12]), .o_data(c_plus_d[136][1]), .i_clk(i_clk));
Add0000000001  u_000000018C_Add0000000001(.i_data_1(matrix_r[393*12+:12]), .i_data_2(matrix_i[393*12+:12]), .o_data(c_plus_d[137][1]), .i_clk(i_clk));
Add0000000001  u_000000018D_Add0000000001(.i_data_1(matrix_r[394*12+:12]), .i_data_2(matrix_i[394*12+:12]), .o_data(c_plus_d[138][1]), .i_clk(i_clk));
Add0000000001  u_000000018E_Add0000000001(.i_data_1(matrix_r[395*12+:12]), .i_data_2(matrix_i[395*12+:12]), .o_data(c_plus_d[139][1]), .i_clk(i_clk));
Add0000000001  u_000000018F_Add0000000001(.i_data_1(matrix_r[396*12+:12]), .i_data_2(matrix_i[396*12+:12]), .o_data(c_plus_d[140][1]), .i_clk(i_clk));
Add0000000001  u_0000000190_Add0000000001(.i_data_1(matrix_r[397*12+:12]), .i_data_2(matrix_i[397*12+:12]), .o_data(c_plus_d[141][1]), .i_clk(i_clk));
Add0000000001  u_0000000191_Add0000000001(.i_data_1(matrix_r[398*12+:12]), .i_data_2(matrix_i[398*12+:12]), .o_data(c_plus_d[142][1]), .i_clk(i_clk));
Add0000000001  u_0000000192_Add0000000001(.i_data_1(matrix_r[399*12+:12]), .i_data_2(matrix_i[399*12+:12]), .o_data(c_plus_d[143][1]), .i_clk(i_clk));
Add0000000001  u_0000000193_Add0000000001(.i_data_1(matrix_r[400*12+:12]), .i_data_2(matrix_i[400*12+:12]), .o_data(c_plus_d[144][1]), .i_clk(i_clk));
Add0000000001  u_0000000194_Add0000000001(.i_data_1(matrix_r[401*12+:12]), .i_data_2(matrix_i[401*12+:12]), .o_data(c_plus_d[145][1]), .i_clk(i_clk));
Add0000000001  u_0000000195_Add0000000001(.i_data_1(matrix_r[402*12+:12]), .i_data_2(matrix_i[402*12+:12]), .o_data(c_plus_d[146][1]), .i_clk(i_clk));
Add0000000001  u_0000000196_Add0000000001(.i_data_1(matrix_r[403*12+:12]), .i_data_2(matrix_i[403*12+:12]), .o_data(c_plus_d[147][1]), .i_clk(i_clk));
Add0000000001  u_0000000197_Add0000000001(.i_data_1(matrix_r[404*12+:12]), .i_data_2(matrix_i[404*12+:12]), .o_data(c_plus_d[148][1]), .i_clk(i_clk));
Add0000000001  u_0000000198_Add0000000001(.i_data_1(matrix_r[405*12+:12]), .i_data_2(matrix_i[405*12+:12]), .o_data(c_plus_d[149][1]), .i_clk(i_clk));
Add0000000001  u_0000000199_Add0000000001(.i_data_1(matrix_r[406*12+:12]), .i_data_2(matrix_i[406*12+:12]), .o_data(c_plus_d[150][1]), .i_clk(i_clk));
Add0000000001  u_000000019A_Add0000000001(.i_data_1(matrix_r[407*12+:12]), .i_data_2(matrix_i[407*12+:12]), .o_data(c_plus_d[151][1]), .i_clk(i_clk));
Add0000000001  u_000000019B_Add0000000001(.i_data_1(matrix_r[408*12+:12]), .i_data_2(matrix_i[408*12+:12]), .o_data(c_plus_d[152][1]), .i_clk(i_clk));
Add0000000001  u_000000019C_Add0000000001(.i_data_1(matrix_r[409*12+:12]), .i_data_2(matrix_i[409*12+:12]), .o_data(c_plus_d[153][1]), .i_clk(i_clk));
Add0000000001  u_000000019D_Add0000000001(.i_data_1(matrix_r[410*12+:12]), .i_data_2(matrix_i[410*12+:12]), .o_data(c_plus_d[154][1]), .i_clk(i_clk));
Add0000000001  u_000000019E_Add0000000001(.i_data_1(matrix_r[411*12+:12]), .i_data_2(matrix_i[411*12+:12]), .o_data(c_plus_d[155][1]), .i_clk(i_clk));
Add0000000001  u_000000019F_Add0000000001(.i_data_1(matrix_r[412*12+:12]), .i_data_2(matrix_i[412*12+:12]), .o_data(c_plus_d[156][1]), .i_clk(i_clk));
Add0000000001  u_00000001A0_Add0000000001(.i_data_1(matrix_r[413*12+:12]), .i_data_2(matrix_i[413*12+:12]), .o_data(c_plus_d[157][1]), .i_clk(i_clk));
Add0000000001  u_00000001A1_Add0000000001(.i_data_1(matrix_r[414*12+:12]), .i_data_2(matrix_i[414*12+:12]), .o_data(c_plus_d[158][1]), .i_clk(i_clk));
Add0000000001  u_00000001A2_Add0000000001(.i_data_1(matrix_r[415*12+:12]), .i_data_2(matrix_i[415*12+:12]), .o_data(c_plus_d[159][1]), .i_clk(i_clk));
Add0000000001  u_00000001A3_Add0000000001(.i_data_1(matrix_r[416*12+:12]), .i_data_2(matrix_i[416*12+:12]), .o_data(c_plus_d[160][1]), .i_clk(i_clk));
Add0000000001  u_00000001A4_Add0000000001(.i_data_1(matrix_r[417*12+:12]), .i_data_2(matrix_i[417*12+:12]), .o_data(c_plus_d[161][1]), .i_clk(i_clk));
Add0000000001  u_00000001A5_Add0000000001(.i_data_1(matrix_r[418*12+:12]), .i_data_2(matrix_i[418*12+:12]), .o_data(c_plus_d[162][1]), .i_clk(i_clk));
Add0000000001  u_00000001A6_Add0000000001(.i_data_1(matrix_r[419*12+:12]), .i_data_2(matrix_i[419*12+:12]), .o_data(c_plus_d[163][1]), .i_clk(i_clk));
Add0000000001  u_00000001A7_Add0000000001(.i_data_1(matrix_r[420*12+:12]), .i_data_2(matrix_i[420*12+:12]), .o_data(c_plus_d[164][1]), .i_clk(i_clk));
Add0000000001  u_00000001A8_Add0000000001(.i_data_1(matrix_r[421*12+:12]), .i_data_2(matrix_i[421*12+:12]), .o_data(c_plus_d[165][1]), .i_clk(i_clk));
Add0000000001  u_00000001A9_Add0000000001(.i_data_1(matrix_r[422*12+:12]), .i_data_2(matrix_i[422*12+:12]), .o_data(c_plus_d[166][1]), .i_clk(i_clk));
Add0000000001  u_00000001AA_Add0000000001(.i_data_1(matrix_r[423*12+:12]), .i_data_2(matrix_i[423*12+:12]), .o_data(c_plus_d[167][1]), .i_clk(i_clk));
Add0000000001  u_00000001AB_Add0000000001(.i_data_1(matrix_r[424*12+:12]), .i_data_2(matrix_i[424*12+:12]), .o_data(c_plus_d[168][1]), .i_clk(i_clk));
Add0000000001  u_00000001AC_Add0000000001(.i_data_1(matrix_r[425*12+:12]), .i_data_2(matrix_i[425*12+:12]), .o_data(c_plus_d[169][1]), .i_clk(i_clk));
Add0000000001  u_00000001AD_Add0000000001(.i_data_1(matrix_r[426*12+:12]), .i_data_2(matrix_i[426*12+:12]), .o_data(c_plus_d[170][1]), .i_clk(i_clk));
Add0000000001  u_00000001AE_Add0000000001(.i_data_1(matrix_r[427*12+:12]), .i_data_2(matrix_i[427*12+:12]), .o_data(c_plus_d[171][1]), .i_clk(i_clk));
Add0000000001  u_00000001AF_Add0000000001(.i_data_1(matrix_r[428*12+:12]), .i_data_2(matrix_i[428*12+:12]), .o_data(c_plus_d[172][1]), .i_clk(i_clk));
Add0000000001  u_00000001B0_Add0000000001(.i_data_1(matrix_r[429*12+:12]), .i_data_2(matrix_i[429*12+:12]), .o_data(c_plus_d[173][1]), .i_clk(i_clk));
Add0000000001  u_00000001B1_Add0000000001(.i_data_1(matrix_r[430*12+:12]), .i_data_2(matrix_i[430*12+:12]), .o_data(c_plus_d[174][1]), .i_clk(i_clk));
Add0000000001  u_00000001B2_Add0000000001(.i_data_1(matrix_r[431*12+:12]), .i_data_2(matrix_i[431*12+:12]), .o_data(c_plus_d[175][1]), .i_clk(i_clk));
Add0000000001  u_00000001B3_Add0000000001(.i_data_1(matrix_r[432*12+:12]), .i_data_2(matrix_i[432*12+:12]), .o_data(c_plus_d[176][1]), .i_clk(i_clk));
Add0000000001  u_00000001B4_Add0000000001(.i_data_1(matrix_r[433*12+:12]), .i_data_2(matrix_i[433*12+:12]), .o_data(c_plus_d[177][1]), .i_clk(i_clk));
Add0000000001  u_00000001B5_Add0000000001(.i_data_1(matrix_r[434*12+:12]), .i_data_2(matrix_i[434*12+:12]), .o_data(c_plus_d[178][1]), .i_clk(i_clk));
Add0000000001  u_00000001B6_Add0000000001(.i_data_1(matrix_r[435*12+:12]), .i_data_2(matrix_i[435*12+:12]), .o_data(c_plus_d[179][1]), .i_clk(i_clk));
Add0000000001  u_00000001B7_Add0000000001(.i_data_1(matrix_r[436*12+:12]), .i_data_2(matrix_i[436*12+:12]), .o_data(c_plus_d[180][1]), .i_clk(i_clk));
Add0000000001  u_00000001B8_Add0000000001(.i_data_1(matrix_r[437*12+:12]), .i_data_2(matrix_i[437*12+:12]), .o_data(c_plus_d[181][1]), .i_clk(i_clk));
Add0000000001  u_00000001B9_Add0000000001(.i_data_1(matrix_r[438*12+:12]), .i_data_2(matrix_i[438*12+:12]), .o_data(c_plus_d[182][1]), .i_clk(i_clk));
Add0000000001  u_00000001BA_Add0000000001(.i_data_1(matrix_r[439*12+:12]), .i_data_2(matrix_i[439*12+:12]), .o_data(c_plus_d[183][1]), .i_clk(i_clk));
Add0000000001  u_00000001BB_Add0000000001(.i_data_1(matrix_r[440*12+:12]), .i_data_2(matrix_i[440*12+:12]), .o_data(c_plus_d[184][1]), .i_clk(i_clk));
Add0000000001  u_00000001BC_Add0000000001(.i_data_1(matrix_r[441*12+:12]), .i_data_2(matrix_i[441*12+:12]), .o_data(c_plus_d[185][1]), .i_clk(i_clk));
Add0000000001  u_00000001BD_Add0000000001(.i_data_1(matrix_r[442*12+:12]), .i_data_2(matrix_i[442*12+:12]), .o_data(c_plus_d[186][1]), .i_clk(i_clk));
Add0000000001  u_00000001BE_Add0000000001(.i_data_1(matrix_r[443*12+:12]), .i_data_2(matrix_i[443*12+:12]), .o_data(c_plus_d[187][1]), .i_clk(i_clk));
Add0000000001  u_00000001BF_Add0000000001(.i_data_1(matrix_r[444*12+:12]), .i_data_2(matrix_i[444*12+:12]), .o_data(c_plus_d[188][1]), .i_clk(i_clk));
Add0000000001  u_00000001C0_Add0000000001(.i_data_1(matrix_r[445*12+:12]), .i_data_2(matrix_i[445*12+:12]), .o_data(c_plus_d[189][1]), .i_clk(i_clk));
Add0000000001  u_00000001C1_Add0000000001(.i_data_1(matrix_r[446*12+:12]), .i_data_2(matrix_i[446*12+:12]), .o_data(c_plus_d[190][1]), .i_clk(i_clk));
Add0000000001  u_00000001C2_Add0000000001(.i_data_1(matrix_r[447*12+:12]), .i_data_2(matrix_i[447*12+:12]), .o_data(c_plus_d[191][1]), .i_clk(i_clk));
Add0000000001  u_00000001C3_Add0000000001(.i_data_1(matrix_r[448*12+:12]), .i_data_2(matrix_i[448*12+:12]), .o_data(c_plus_d[192][1]), .i_clk(i_clk));
Add0000000001  u_00000001C4_Add0000000001(.i_data_1(matrix_r[449*12+:12]), .i_data_2(matrix_i[449*12+:12]), .o_data(c_plus_d[193][1]), .i_clk(i_clk));
Add0000000001  u_00000001C5_Add0000000001(.i_data_1(matrix_r[450*12+:12]), .i_data_2(matrix_i[450*12+:12]), .o_data(c_plus_d[194][1]), .i_clk(i_clk));
Add0000000001  u_00000001C6_Add0000000001(.i_data_1(matrix_r[451*12+:12]), .i_data_2(matrix_i[451*12+:12]), .o_data(c_plus_d[195][1]), .i_clk(i_clk));
Add0000000001  u_00000001C7_Add0000000001(.i_data_1(matrix_r[452*12+:12]), .i_data_2(matrix_i[452*12+:12]), .o_data(c_plus_d[196][1]), .i_clk(i_clk));
Add0000000001  u_00000001C8_Add0000000001(.i_data_1(matrix_r[453*12+:12]), .i_data_2(matrix_i[453*12+:12]), .o_data(c_plus_d[197][1]), .i_clk(i_clk));
Add0000000001  u_00000001C9_Add0000000001(.i_data_1(matrix_r[454*12+:12]), .i_data_2(matrix_i[454*12+:12]), .o_data(c_plus_d[198][1]), .i_clk(i_clk));
Add0000000001  u_00000001CA_Add0000000001(.i_data_1(matrix_r[455*12+:12]), .i_data_2(matrix_i[455*12+:12]), .o_data(c_plus_d[199][1]), .i_clk(i_clk));
Add0000000001  u_00000001CB_Add0000000001(.i_data_1(matrix_r[456*12+:12]), .i_data_2(matrix_i[456*12+:12]), .o_data(c_plus_d[200][1]), .i_clk(i_clk));
Add0000000001  u_00000001CC_Add0000000001(.i_data_1(matrix_r[457*12+:12]), .i_data_2(matrix_i[457*12+:12]), .o_data(c_plus_d[201][1]), .i_clk(i_clk));
Add0000000001  u_00000001CD_Add0000000001(.i_data_1(matrix_r[458*12+:12]), .i_data_2(matrix_i[458*12+:12]), .o_data(c_plus_d[202][1]), .i_clk(i_clk));
Add0000000001  u_00000001CE_Add0000000001(.i_data_1(matrix_r[459*12+:12]), .i_data_2(matrix_i[459*12+:12]), .o_data(c_plus_d[203][1]), .i_clk(i_clk));
Add0000000001  u_00000001CF_Add0000000001(.i_data_1(matrix_r[460*12+:12]), .i_data_2(matrix_i[460*12+:12]), .o_data(c_plus_d[204][1]), .i_clk(i_clk));
Add0000000001  u_00000001D0_Add0000000001(.i_data_1(matrix_r[461*12+:12]), .i_data_2(matrix_i[461*12+:12]), .o_data(c_plus_d[205][1]), .i_clk(i_clk));
Add0000000001  u_00000001D1_Add0000000001(.i_data_1(matrix_r[462*12+:12]), .i_data_2(matrix_i[462*12+:12]), .o_data(c_plus_d[206][1]), .i_clk(i_clk));
Add0000000001  u_00000001D2_Add0000000001(.i_data_1(matrix_r[463*12+:12]), .i_data_2(matrix_i[463*12+:12]), .o_data(c_plus_d[207][1]), .i_clk(i_clk));
Add0000000001  u_00000001D3_Add0000000001(.i_data_1(matrix_r[464*12+:12]), .i_data_2(matrix_i[464*12+:12]), .o_data(c_plus_d[208][1]), .i_clk(i_clk));
Add0000000001  u_00000001D4_Add0000000001(.i_data_1(matrix_r[465*12+:12]), .i_data_2(matrix_i[465*12+:12]), .o_data(c_plus_d[209][1]), .i_clk(i_clk));
Add0000000001  u_00000001D5_Add0000000001(.i_data_1(matrix_r[466*12+:12]), .i_data_2(matrix_i[466*12+:12]), .o_data(c_plus_d[210][1]), .i_clk(i_clk));
Add0000000001  u_00000001D6_Add0000000001(.i_data_1(matrix_r[467*12+:12]), .i_data_2(matrix_i[467*12+:12]), .o_data(c_plus_d[211][1]), .i_clk(i_clk));
Add0000000001  u_00000001D7_Add0000000001(.i_data_1(matrix_r[468*12+:12]), .i_data_2(matrix_i[468*12+:12]), .o_data(c_plus_d[212][1]), .i_clk(i_clk));
Add0000000001  u_00000001D8_Add0000000001(.i_data_1(matrix_r[469*12+:12]), .i_data_2(matrix_i[469*12+:12]), .o_data(c_plus_d[213][1]), .i_clk(i_clk));
Add0000000001  u_00000001D9_Add0000000001(.i_data_1(matrix_r[470*12+:12]), .i_data_2(matrix_i[470*12+:12]), .o_data(c_plus_d[214][1]), .i_clk(i_clk));
Add0000000001  u_00000001DA_Add0000000001(.i_data_1(matrix_r[471*12+:12]), .i_data_2(matrix_i[471*12+:12]), .o_data(c_plus_d[215][1]), .i_clk(i_clk));
Add0000000001  u_00000001DB_Add0000000001(.i_data_1(matrix_r[472*12+:12]), .i_data_2(matrix_i[472*12+:12]), .o_data(c_plus_d[216][1]), .i_clk(i_clk));
Add0000000001  u_00000001DC_Add0000000001(.i_data_1(matrix_r[473*12+:12]), .i_data_2(matrix_i[473*12+:12]), .o_data(c_plus_d[217][1]), .i_clk(i_clk));
Add0000000001  u_00000001DD_Add0000000001(.i_data_1(matrix_r[474*12+:12]), .i_data_2(matrix_i[474*12+:12]), .o_data(c_plus_d[218][1]), .i_clk(i_clk));
Add0000000001  u_00000001DE_Add0000000001(.i_data_1(matrix_r[475*12+:12]), .i_data_2(matrix_i[475*12+:12]), .o_data(c_plus_d[219][1]), .i_clk(i_clk));
Add0000000001  u_00000001DF_Add0000000001(.i_data_1(matrix_r[476*12+:12]), .i_data_2(matrix_i[476*12+:12]), .o_data(c_plus_d[220][1]), .i_clk(i_clk));
Add0000000001  u_00000001E0_Add0000000001(.i_data_1(matrix_r[477*12+:12]), .i_data_2(matrix_i[477*12+:12]), .o_data(c_plus_d[221][1]), .i_clk(i_clk));
Add0000000001  u_00000001E1_Add0000000001(.i_data_1(matrix_r[478*12+:12]), .i_data_2(matrix_i[478*12+:12]), .o_data(c_plus_d[222][1]), .i_clk(i_clk));
Add0000000001  u_00000001E2_Add0000000001(.i_data_1(matrix_r[479*12+:12]), .i_data_2(matrix_i[479*12+:12]), .o_data(c_plus_d[223][1]), .i_clk(i_clk));
Add0000000001  u_00000001E3_Add0000000001(.i_data_1(matrix_r[480*12+:12]), .i_data_2(matrix_i[480*12+:12]), .o_data(c_plus_d[224][1]), .i_clk(i_clk));
Add0000000001  u_00000001E4_Add0000000001(.i_data_1(matrix_r[481*12+:12]), .i_data_2(matrix_i[481*12+:12]), .o_data(c_plus_d[225][1]), .i_clk(i_clk));
Add0000000001  u_00000001E5_Add0000000001(.i_data_1(matrix_r[482*12+:12]), .i_data_2(matrix_i[482*12+:12]), .o_data(c_plus_d[226][1]), .i_clk(i_clk));
Add0000000001  u_00000001E6_Add0000000001(.i_data_1(matrix_r[483*12+:12]), .i_data_2(matrix_i[483*12+:12]), .o_data(c_plus_d[227][1]), .i_clk(i_clk));
Add0000000001  u_00000001E7_Add0000000001(.i_data_1(matrix_r[484*12+:12]), .i_data_2(matrix_i[484*12+:12]), .o_data(c_plus_d[228][1]), .i_clk(i_clk));
Add0000000001  u_00000001E8_Add0000000001(.i_data_1(matrix_r[485*12+:12]), .i_data_2(matrix_i[485*12+:12]), .o_data(c_plus_d[229][1]), .i_clk(i_clk));
Add0000000001  u_00000001E9_Add0000000001(.i_data_1(matrix_r[486*12+:12]), .i_data_2(matrix_i[486*12+:12]), .o_data(c_plus_d[230][1]), .i_clk(i_clk));
Add0000000001  u_00000001EA_Add0000000001(.i_data_1(matrix_r[487*12+:12]), .i_data_2(matrix_i[487*12+:12]), .o_data(c_plus_d[231][1]), .i_clk(i_clk));
Add0000000001  u_00000001EB_Add0000000001(.i_data_1(matrix_r[488*12+:12]), .i_data_2(matrix_i[488*12+:12]), .o_data(c_plus_d[232][1]), .i_clk(i_clk));
Add0000000001  u_00000001EC_Add0000000001(.i_data_1(matrix_r[489*12+:12]), .i_data_2(matrix_i[489*12+:12]), .o_data(c_plus_d[233][1]), .i_clk(i_clk));
Add0000000001  u_00000001ED_Add0000000001(.i_data_1(matrix_r[490*12+:12]), .i_data_2(matrix_i[490*12+:12]), .o_data(c_plus_d[234][1]), .i_clk(i_clk));
Add0000000001  u_00000001EE_Add0000000001(.i_data_1(matrix_r[491*12+:12]), .i_data_2(matrix_i[491*12+:12]), .o_data(c_plus_d[235][1]), .i_clk(i_clk));
Add0000000001  u_00000001EF_Add0000000001(.i_data_1(matrix_r[492*12+:12]), .i_data_2(matrix_i[492*12+:12]), .o_data(c_plus_d[236][1]), .i_clk(i_clk));
Add0000000001  u_00000001F0_Add0000000001(.i_data_1(matrix_r[493*12+:12]), .i_data_2(matrix_i[493*12+:12]), .o_data(c_plus_d[237][1]), .i_clk(i_clk));
Add0000000001  u_00000001F1_Add0000000001(.i_data_1(matrix_r[494*12+:12]), .i_data_2(matrix_i[494*12+:12]), .o_data(c_plus_d[238][1]), .i_clk(i_clk));
Add0000000001  u_00000001F2_Add0000000001(.i_data_1(matrix_r[495*12+:12]), .i_data_2(matrix_i[495*12+:12]), .o_data(c_plus_d[239][1]), .i_clk(i_clk));
Add0000000001  u_00000001F3_Add0000000001(.i_data_1(matrix_r[496*12+:12]), .i_data_2(matrix_i[496*12+:12]), .o_data(c_plus_d[240][1]), .i_clk(i_clk));
Add0000000001  u_00000001F4_Add0000000001(.i_data_1(matrix_r[497*12+:12]), .i_data_2(matrix_i[497*12+:12]), .o_data(c_plus_d[241][1]), .i_clk(i_clk));
Add0000000001  u_00000001F5_Add0000000001(.i_data_1(matrix_r[498*12+:12]), .i_data_2(matrix_i[498*12+:12]), .o_data(c_plus_d[242][1]), .i_clk(i_clk));
Add0000000001  u_00000001F6_Add0000000001(.i_data_1(matrix_r[499*12+:12]), .i_data_2(matrix_i[499*12+:12]), .o_data(c_plus_d[243][1]), .i_clk(i_clk));
Add0000000001  u_00000001F7_Add0000000001(.i_data_1(matrix_r[500*12+:12]), .i_data_2(matrix_i[500*12+:12]), .o_data(c_plus_d[244][1]), .i_clk(i_clk));
Add0000000001  u_00000001F8_Add0000000001(.i_data_1(matrix_r[501*12+:12]), .i_data_2(matrix_i[501*12+:12]), .o_data(c_plus_d[245][1]), .i_clk(i_clk));
Add0000000001  u_00000001F9_Add0000000001(.i_data_1(matrix_r[502*12+:12]), .i_data_2(matrix_i[502*12+:12]), .o_data(c_plus_d[246][1]), .i_clk(i_clk));
Add0000000001  u_00000001FA_Add0000000001(.i_data_1(matrix_r[503*12+:12]), .i_data_2(matrix_i[503*12+:12]), .o_data(c_plus_d[247][1]), .i_clk(i_clk));
Add0000000001  u_00000001FB_Add0000000001(.i_data_1(matrix_r[504*12+:12]), .i_data_2(matrix_i[504*12+:12]), .o_data(c_plus_d[248][1]), .i_clk(i_clk));
Add0000000001  u_00000001FC_Add0000000001(.i_data_1(matrix_r[505*12+:12]), .i_data_2(matrix_i[505*12+:12]), .o_data(c_plus_d[249][1]), .i_clk(i_clk));
Add0000000001  u_00000001FD_Add0000000001(.i_data_1(matrix_r[506*12+:12]), .i_data_2(matrix_i[506*12+:12]), .o_data(c_plus_d[250][1]), .i_clk(i_clk));
Add0000000001  u_00000001FE_Add0000000001(.i_data_1(matrix_r[507*12+:12]), .i_data_2(matrix_i[507*12+:12]), .o_data(c_plus_d[251][1]), .i_clk(i_clk));
Add0000000001  u_00000001FF_Add0000000001(.i_data_1(matrix_r[508*12+:12]), .i_data_2(matrix_i[508*12+:12]), .o_data(c_plus_d[252][1]), .i_clk(i_clk));
Add0000000001  u_0000000200_Add0000000001(.i_data_1(matrix_r[509*12+:12]), .i_data_2(matrix_i[509*12+:12]), .o_data(c_plus_d[253][1]), .i_clk(i_clk));
Add0000000001  u_0000000201_Add0000000001(.i_data_1(matrix_r[510*12+:12]), .i_data_2(matrix_i[510*12+:12]), .o_data(c_plus_d[254][1]), .i_clk(i_clk));
Add0000000001  u_0000000202_Add0000000001(.i_data_1(matrix_r[511*12+:12]), .i_data_2(matrix_i[511*12+:12]), .o_data(c_plus_d[255][1]), .i_clk(i_clk));
Add0000000001  u_0000000203_Add0000000001(.i_data_1(vector_r[2*12+:12]), .i_data_2(vector_i[2*12+:12]), .o_data(a_plus_b[2]), .i_clk(i_clk));
Sub0000000001  u_0000000003_Sub0000000001(.i_data_1(vector_i[2*12+:12]), .i_data_2(vector_r[2*12+:12]), .o_data(b_minus_a[2]), .i_clk(i_clk));
Add0000000001  u_0000000204_Add0000000001(.i_data_1(matrix_r[512*12+:12]), .i_data_2(matrix_i[512*12+:12]), .o_data(c_plus_d[0][2]), .i_clk(i_clk));
Add0000000001  u_0000000205_Add0000000001(.i_data_1(matrix_r[513*12+:12]), .i_data_2(matrix_i[513*12+:12]), .o_data(c_plus_d[1][2]), .i_clk(i_clk));
Add0000000001  u_0000000206_Add0000000001(.i_data_1(matrix_r[514*12+:12]), .i_data_2(matrix_i[514*12+:12]), .o_data(c_plus_d[2][2]), .i_clk(i_clk));
Add0000000001  u_0000000207_Add0000000001(.i_data_1(matrix_r[515*12+:12]), .i_data_2(matrix_i[515*12+:12]), .o_data(c_plus_d[3][2]), .i_clk(i_clk));
Add0000000001  u_0000000208_Add0000000001(.i_data_1(matrix_r[516*12+:12]), .i_data_2(matrix_i[516*12+:12]), .o_data(c_plus_d[4][2]), .i_clk(i_clk));
Add0000000001  u_0000000209_Add0000000001(.i_data_1(matrix_r[517*12+:12]), .i_data_2(matrix_i[517*12+:12]), .o_data(c_plus_d[5][2]), .i_clk(i_clk));
Add0000000001  u_000000020A_Add0000000001(.i_data_1(matrix_r[518*12+:12]), .i_data_2(matrix_i[518*12+:12]), .o_data(c_plus_d[6][2]), .i_clk(i_clk));
Add0000000001  u_000000020B_Add0000000001(.i_data_1(matrix_r[519*12+:12]), .i_data_2(matrix_i[519*12+:12]), .o_data(c_plus_d[7][2]), .i_clk(i_clk));
Add0000000001  u_000000020C_Add0000000001(.i_data_1(matrix_r[520*12+:12]), .i_data_2(matrix_i[520*12+:12]), .o_data(c_plus_d[8][2]), .i_clk(i_clk));
Add0000000001  u_000000020D_Add0000000001(.i_data_1(matrix_r[521*12+:12]), .i_data_2(matrix_i[521*12+:12]), .o_data(c_plus_d[9][2]), .i_clk(i_clk));
Add0000000001  u_000000020E_Add0000000001(.i_data_1(matrix_r[522*12+:12]), .i_data_2(matrix_i[522*12+:12]), .o_data(c_plus_d[10][2]), .i_clk(i_clk));
Add0000000001  u_000000020F_Add0000000001(.i_data_1(matrix_r[523*12+:12]), .i_data_2(matrix_i[523*12+:12]), .o_data(c_plus_d[11][2]), .i_clk(i_clk));
Add0000000001  u_0000000210_Add0000000001(.i_data_1(matrix_r[524*12+:12]), .i_data_2(matrix_i[524*12+:12]), .o_data(c_plus_d[12][2]), .i_clk(i_clk));
Add0000000001  u_0000000211_Add0000000001(.i_data_1(matrix_r[525*12+:12]), .i_data_2(matrix_i[525*12+:12]), .o_data(c_plus_d[13][2]), .i_clk(i_clk));
Add0000000001  u_0000000212_Add0000000001(.i_data_1(matrix_r[526*12+:12]), .i_data_2(matrix_i[526*12+:12]), .o_data(c_plus_d[14][2]), .i_clk(i_clk));
Add0000000001  u_0000000213_Add0000000001(.i_data_1(matrix_r[527*12+:12]), .i_data_2(matrix_i[527*12+:12]), .o_data(c_plus_d[15][2]), .i_clk(i_clk));
Add0000000001  u_0000000214_Add0000000001(.i_data_1(matrix_r[528*12+:12]), .i_data_2(matrix_i[528*12+:12]), .o_data(c_plus_d[16][2]), .i_clk(i_clk));
Add0000000001  u_0000000215_Add0000000001(.i_data_1(matrix_r[529*12+:12]), .i_data_2(matrix_i[529*12+:12]), .o_data(c_plus_d[17][2]), .i_clk(i_clk));
Add0000000001  u_0000000216_Add0000000001(.i_data_1(matrix_r[530*12+:12]), .i_data_2(matrix_i[530*12+:12]), .o_data(c_plus_d[18][2]), .i_clk(i_clk));
Add0000000001  u_0000000217_Add0000000001(.i_data_1(matrix_r[531*12+:12]), .i_data_2(matrix_i[531*12+:12]), .o_data(c_plus_d[19][2]), .i_clk(i_clk));
Add0000000001  u_0000000218_Add0000000001(.i_data_1(matrix_r[532*12+:12]), .i_data_2(matrix_i[532*12+:12]), .o_data(c_plus_d[20][2]), .i_clk(i_clk));
Add0000000001  u_0000000219_Add0000000001(.i_data_1(matrix_r[533*12+:12]), .i_data_2(matrix_i[533*12+:12]), .o_data(c_plus_d[21][2]), .i_clk(i_clk));
Add0000000001  u_000000021A_Add0000000001(.i_data_1(matrix_r[534*12+:12]), .i_data_2(matrix_i[534*12+:12]), .o_data(c_plus_d[22][2]), .i_clk(i_clk));
Add0000000001  u_000000021B_Add0000000001(.i_data_1(matrix_r[535*12+:12]), .i_data_2(matrix_i[535*12+:12]), .o_data(c_plus_d[23][2]), .i_clk(i_clk));
Add0000000001  u_000000021C_Add0000000001(.i_data_1(matrix_r[536*12+:12]), .i_data_2(matrix_i[536*12+:12]), .o_data(c_plus_d[24][2]), .i_clk(i_clk));
Add0000000001  u_000000021D_Add0000000001(.i_data_1(matrix_r[537*12+:12]), .i_data_2(matrix_i[537*12+:12]), .o_data(c_plus_d[25][2]), .i_clk(i_clk));
Add0000000001  u_000000021E_Add0000000001(.i_data_1(matrix_r[538*12+:12]), .i_data_2(matrix_i[538*12+:12]), .o_data(c_plus_d[26][2]), .i_clk(i_clk));
Add0000000001  u_000000021F_Add0000000001(.i_data_1(matrix_r[539*12+:12]), .i_data_2(matrix_i[539*12+:12]), .o_data(c_plus_d[27][2]), .i_clk(i_clk));
Add0000000001  u_0000000220_Add0000000001(.i_data_1(matrix_r[540*12+:12]), .i_data_2(matrix_i[540*12+:12]), .o_data(c_plus_d[28][2]), .i_clk(i_clk));
Add0000000001  u_0000000221_Add0000000001(.i_data_1(matrix_r[541*12+:12]), .i_data_2(matrix_i[541*12+:12]), .o_data(c_plus_d[29][2]), .i_clk(i_clk));
Add0000000001  u_0000000222_Add0000000001(.i_data_1(matrix_r[542*12+:12]), .i_data_2(matrix_i[542*12+:12]), .o_data(c_plus_d[30][2]), .i_clk(i_clk));
Add0000000001  u_0000000223_Add0000000001(.i_data_1(matrix_r[543*12+:12]), .i_data_2(matrix_i[543*12+:12]), .o_data(c_plus_d[31][2]), .i_clk(i_clk));
Add0000000001  u_0000000224_Add0000000001(.i_data_1(matrix_r[544*12+:12]), .i_data_2(matrix_i[544*12+:12]), .o_data(c_plus_d[32][2]), .i_clk(i_clk));
Add0000000001  u_0000000225_Add0000000001(.i_data_1(matrix_r[545*12+:12]), .i_data_2(matrix_i[545*12+:12]), .o_data(c_plus_d[33][2]), .i_clk(i_clk));
Add0000000001  u_0000000226_Add0000000001(.i_data_1(matrix_r[546*12+:12]), .i_data_2(matrix_i[546*12+:12]), .o_data(c_plus_d[34][2]), .i_clk(i_clk));
Add0000000001  u_0000000227_Add0000000001(.i_data_1(matrix_r[547*12+:12]), .i_data_2(matrix_i[547*12+:12]), .o_data(c_plus_d[35][2]), .i_clk(i_clk));
Add0000000001  u_0000000228_Add0000000001(.i_data_1(matrix_r[548*12+:12]), .i_data_2(matrix_i[548*12+:12]), .o_data(c_plus_d[36][2]), .i_clk(i_clk));
Add0000000001  u_0000000229_Add0000000001(.i_data_1(matrix_r[549*12+:12]), .i_data_2(matrix_i[549*12+:12]), .o_data(c_plus_d[37][2]), .i_clk(i_clk));
Add0000000001  u_000000022A_Add0000000001(.i_data_1(matrix_r[550*12+:12]), .i_data_2(matrix_i[550*12+:12]), .o_data(c_plus_d[38][2]), .i_clk(i_clk));
Add0000000001  u_000000022B_Add0000000001(.i_data_1(matrix_r[551*12+:12]), .i_data_2(matrix_i[551*12+:12]), .o_data(c_plus_d[39][2]), .i_clk(i_clk));
Add0000000001  u_000000022C_Add0000000001(.i_data_1(matrix_r[552*12+:12]), .i_data_2(matrix_i[552*12+:12]), .o_data(c_plus_d[40][2]), .i_clk(i_clk));
Add0000000001  u_000000022D_Add0000000001(.i_data_1(matrix_r[553*12+:12]), .i_data_2(matrix_i[553*12+:12]), .o_data(c_plus_d[41][2]), .i_clk(i_clk));
Add0000000001  u_000000022E_Add0000000001(.i_data_1(matrix_r[554*12+:12]), .i_data_2(matrix_i[554*12+:12]), .o_data(c_plus_d[42][2]), .i_clk(i_clk));
Add0000000001  u_000000022F_Add0000000001(.i_data_1(matrix_r[555*12+:12]), .i_data_2(matrix_i[555*12+:12]), .o_data(c_plus_d[43][2]), .i_clk(i_clk));
Add0000000001  u_0000000230_Add0000000001(.i_data_1(matrix_r[556*12+:12]), .i_data_2(matrix_i[556*12+:12]), .o_data(c_plus_d[44][2]), .i_clk(i_clk));
Add0000000001  u_0000000231_Add0000000001(.i_data_1(matrix_r[557*12+:12]), .i_data_2(matrix_i[557*12+:12]), .o_data(c_plus_d[45][2]), .i_clk(i_clk));
Add0000000001  u_0000000232_Add0000000001(.i_data_1(matrix_r[558*12+:12]), .i_data_2(matrix_i[558*12+:12]), .o_data(c_plus_d[46][2]), .i_clk(i_clk));
Add0000000001  u_0000000233_Add0000000001(.i_data_1(matrix_r[559*12+:12]), .i_data_2(matrix_i[559*12+:12]), .o_data(c_plus_d[47][2]), .i_clk(i_clk));
Add0000000001  u_0000000234_Add0000000001(.i_data_1(matrix_r[560*12+:12]), .i_data_2(matrix_i[560*12+:12]), .o_data(c_plus_d[48][2]), .i_clk(i_clk));
Add0000000001  u_0000000235_Add0000000001(.i_data_1(matrix_r[561*12+:12]), .i_data_2(matrix_i[561*12+:12]), .o_data(c_plus_d[49][2]), .i_clk(i_clk));
Add0000000001  u_0000000236_Add0000000001(.i_data_1(matrix_r[562*12+:12]), .i_data_2(matrix_i[562*12+:12]), .o_data(c_plus_d[50][2]), .i_clk(i_clk));
Add0000000001  u_0000000237_Add0000000001(.i_data_1(matrix_r[563*12+:12]), .i_data_2(matrix_i[563*12+:12]), .o_data(c_plus_d[51][2]), .i_clk(i_clk));
Add0000000001  u_0000000238_Add0000000001(.i_data_1(matrix_r[564*12+:12]), .i_data_2(matrix_i[564*12+:12]), .o_data(c_plus_d[52][2]), .i_clk(i_clk));
Add0000000001  u_0000000239_Add0000000001(.i_data_1(matrix_r[565*12+:12]), .i_data_2(matrix_i[565*12+:12]), .o_data(c_plus_d[53][2]), .i_clk(i_clk));
Add0000000001  u_000000023A_Add0000000001(.i_data_1(matrix_r[566*12+:12]), .i_data_2(matrix_i[566*12+:12]), .o_data(c_plus_d[54][2]), .i_clk(i_clk));
Add0000000001  u_000000023B_Add0000000001(.i_data_1(matrix_r[567*12+:12]), .i_data_2(matrix_i[567*12+:12]), .o_data(c_plus_d[55][2]), .i_clk(i_clk));
Add0000000001  u_000000023C_Add0000000001(.i_data_1(matrix_r[568*12+:12]), .i_data_2(matrix_i[568*12+:12]), .o_data(c_plus_d[56][2]), .i_clk(i_clk));
Add0000000001  u_000000023D_Add0000000001(.i_data_1(matrix_r[569*12+:12]), .i_data_2(matrix_i[569*12+:12]), .o_data(c_plus_d[57][2]), .i_clk(i_clk));
Add0000000001  u_000000023E_Add0000000001(.i_data_1(matrix_r[570*12+:12]), .i_data_2(matrix_i[570*12+:12]), .o_data(c_plus_d[58][2]), .i_clk(i_clk));
Add0000000001  u_000000023F_Add0000000001(.i_data_1(matrix_r[571*12+:12]), .i_data_2(matrix_i[571*12+:12]), .o_data(c_plus_d[59][2]), .i_clk(i_clk));
Add0000000001  u_0000000240_Add0000000001(.i_data_1(matrix_r[572*12+:12]), .i_data_2(matrix_i[572*12+:12]), .o_data(c_plus_d[60][2]), .i_clk(i_clk));
Add0000000001  u_0000000241_Add0000000001(.i_data_1(matrix_r[573*12+:12]), .i_data_2(matrix_i[573*12+:12]), .o_data(c_plus_d[61][2]), .i_clk(i_clk));
Add0000000001  u_0000000242_Add0000000001(.i_data_1(matrix_r[574*12+:12]), .i_data_2(matrix_i[574*12+:12]), .o_data(c_plus_d[62][2]), .i_clk(i_clk));
Add0000000001  u_0000000243_Add0000000001(.i_data_1(matrix_r[575*12+:12]), .i_data_2(matrix_i[575*12+:12]), .o_data(c_plus_d[63][2]), .i_clk(i_clk));
Add0000000001  u_0000000244_Add0000000001(.i_data_1(matrix_r[576*12+:12]), .i_data_2(matrix_i[576*12+:12]), .o_data(c_plus_d[64][2]), .i_clk(i_clk));
Add0000000001  u_0000000245_Add0000000001(.i_data_1(matrix_r[577*12+:12]), .i_data_2(matrix_i[577*12+:12]), .o_data(c_plus_d[65][2]), .i_clk(i_clk));
Add0000000001  u_0000000246_Add0000000001(.i_data_1(matrix_r[578*12+:12]), .i_data_2(matrix_i[578*12+:12]), .o_data(c_plus_d[66][2]), .i_clk(i_clk));
Add0000000001  u_0000000247_Add0000000001(.i_data_1(matrix_r[579*12+:12]), .i_data_2(matrix_i[579*12+:12]), .o_data(c_plus_d[67][2]), .i_clk(i_clk));
Add0000000001  u_0000000248_Add0000000001(.i_data_1(matrix_r[580*12+:12]), .i_data_2(matrix_i[580*12+:12]), .o_data(c_plus_d[68][2]), .i_clk(i_clk));
Add0000000001  u_0000000249_Add0000000001(.i_data_1(matrix_r[581*12+:12]), .i_data_2(matrix_i[581*12+:12]), .o_data(c_plus_d[69][2]), .i_clk(i_clk));
Add0000000001  u_000000024A_Add0000000001(.i_data_1(matrix_r[582*12+:12]), .i_data_2(matrix_i[582*12+:12]), .o_data(c_plus_d[70][2]), .i_clk(i_clk));
Add0000000001  u_000000024B_Add0000000001(.i_data_1(matrix_r[583*12+:12]), .i_data_2(matrix_i[583*12+:12]), .o_data(c_plus_d[71][2]), .i_clk(i_clk));
Add0000000001  u_000000024C_Add0000000001(.i_data_1(matrix_r[584*12+:12]), .i_data_2(matrix_i[584*12+:12]), .o_data(c_plus_d[72][2]), .i_clk(i_clk));
Add0000000001  u_000000024D_Add0000000001(.i_data_1(matrix_r[585*12+:12]), .i_data_2(matrix_i[585*12+:12]), .o_data(c_plus_d[73][2]), .i_clk(i_clk));
Add0000000001  u_000000024E_Add0000000001(.i_data_1(matrix_r[586*12+:12]), .i_data_2(matrix_i[586*12+:12]), .o_data(c_plus_d[74][2]), .i_clk(i_clk));
Add0000000001  u_000000024F_Add0000000001(.i_data_1(matrix_r[587*12+:12]), .i_data_2(matrix_i[587*12+:12]), .o_data(c_plus_d[75][2]), .i_clk(i_clk));
Add0000000001  u_0000000250_Add0000000001(.i_data_1(matrix_r[588*12+:12]), .i_data_2(matrix_i[588*12+:12]), .o_data(c_plus_d[76][2]), .i_clk(i_clk));
Add0000000001  u_0000000251_Add0000000001(.i_data_1(matrix_r[589*12+:12]), .i_data_2(matrix_i[589*12+:12]), .o_data(c_plus_d[77][2]), .i_clk(i_clk));
Add0000000001  u_0000000252_Add0000000001(.i_data_1(matrix_r[590*12+:12]), .i_data_2(matrix_i[590*12+:12]), .o_data(c_plus_d[78][2]), .i_clk(i_clk));
Add0000000001  u_0000000253_Add0000000001(.i_data_1(matrix_r[591*12+:12]), .i_data_2(matrix_i[591*12+:12]), .o_data(c_plus_d[79][2]), .i_clk(i_clk));
Add0000000001  u_0000000254_Add0000000001(.i_data_1(matrix_r[592*12+:12]), .i_data_2(matrix_i[592*12+:12]), .o_data(c_plus_d[80][2]), .i_clk(i_clk));
Add0000000001  u_0000000255_Add0000000001(.i_data_1(matrix_r[593*12+:12]), .i_data_2(matrix_i[593*12+:12]), .o_data(c_plus_d[81][2]), .i_clk(i_clk));
Add0000000001  u_0000000256_Add0000000001(.i_data_1(matrix_r[594*12+:12]), .i_data_2(matrix_i[594*12+:12]), .o_data(c_plus_d[82][2]), .i_clk(i_clk));
Add0000000001  u_0000000257_Add0000000001(.i_data_1(matrix_r[595*12+:12]), .i_data_2(matrix_i[595*12+:12]), .o_data(c_plus_d[83][2]), .i_clk(i_clk));
Add0000000001  u_0000000258_Add0000000001(.i_data_1(matrix_r[596*12+:12]), .i_data_2(matrix_i[596*12+:12]), .o_data(c_plus_d[84][2]), .i_clk(i_clk));
Add0000000001  u_0000000259_Add0000000001(.i_data_1(matrix_r[597*12+:12]), .i_data_2(matrix_i[597*12+:12]), .o_data(c_plus_d[85][2]), .i_clk(i_clk));
Add0000000001  u_000000025A_Add0000000001(.i_data_1(matrix_r[598*12+:12]), .i_data_2(matrix_i[598*12+:12]), .o_data(c_plus_d[86][2]), .i_clk(i_clk));
Add0000000001  u_000000025B_Add0000000001(.i_data_1(matrix_r[599*12+:12]), .i_data_2(matrix_i[599*12+:12]), .o_data(c_plus_d[87][2]), .i_clk(i_clk));
Add0000000001  u_000000025C_Add0000000001(.i_data_1(matrix_r[600*12+:12]), .i_data_2(matrix_i[600*12+:12]), .o_data(c_plus_d[88][2]), .i_clk(i_clk));
Add0000000001  u_000000025D_Add0000000001(.i_data_1(matrix_r[601*12+:12]), .i_data_2(matrix_i[601*12+:12]), .o_data(c_plus_d[89][2]), .i_clk(i_clk));
Add0000000001  u_000000025E_Add0000000001(.i_data_1(matrix_r[602*12+:12]), .i_data_2(matrix_i[602*12+:12]), .o_data(c_plus_d[90][2]), .i_clk(i_clk));
Add0000000001  u_000000025F_Add0000000001(.i_data_1(matrix_r[603*12+:12]), .i_data_2(matrix_i[603*12+:12]), .o_data(c_plus_d[91][2]), .i_clk(i_clk));
Add0000000001  u_0000000260_Add0000000001(.i_data_1(matrix_r[604*12+:12]), .i_data_2(matrix_i[604*12+:12]), .o_data(c_plus_d[92][2]), .i_clk(i_clk));
Add0000000001  u_0000000261_Add0000000001(.i_data_1(matrix_r[605*12+:12]), .i_data_2(matrix_i[605*12+:12]), .o_data(c_plus_d[93][2]), .i_clk(i_clk));
Add0000000001  u_0000000262_Add0000000001(.i_data_1(matrix_r[606*12+:12]), .i_data_2(matrix_i[606*12+:12]), .o_data(c_plus_d[94][2]), .i_clk(i_clk));
Add0000000001  u_0000000263_Add0000000001(.i_data_1(matrix_r[607*12+:12]), .i_data_2(matrix_i[607*12+:12]), .o_data(c_plus_d[95][2]), .i_clk(i_clk));
Add0000000001  u_0000000264_Add0000000001(.i_data_1(matrix_r[608*12+:12]), .i_data_2(matrix_i[608*12+:12]), .o_data(c_plus_d[96][2]), .i_clk(i_clk));
Add0000000001  u_0000000265_Add0000000001(.i_data_1(matrix_r[609*12+:12]), .i_data_2(matrix_i[609*12+:12]), .o_data(c_plus_d[97][2]), .i_clk(i_clk));
Add0000000001  u_0000000266_Add0000000001(.i_data_1(matrix_r[610*12+:12]), .i_data_2(matrix_i[610*12+:12]), .o_data(c_plus_d[98][2]), .i_clk(i_clk));
Add0000000001  u_0000000267_Add0000000001(.i_data_1(matrix_r[611*12+:12]), .i_data_2(matrix_i[611*12+:12]), .o_data(c_plus_d[99][2]), .i_clk(i_clk));
Add0000000001  u_0000000268_Add0000000001(.i_data_1(matrix_r[612*12+:12]), .i_data_2(matrix_i[612*12+:12]), .o_data(c_plus_d[100][2]), .i_clk(i_clk));
Add0000000001  u_0000000269_Add0000000001(.i_data_1(matrix_r[613*12+:12]), .i_data_2(matrix_i[613*12+:12]), .o_data(c_plus_d[101][2]), .i_clk(i_clk));
Add0000000001  u_000000026A_Add0000000001(.i_data_1(matrix_r[614*12+:12]), .i_data_2(matrix_i[614*12+:12]), .o_data(c_plus_d[102][2]), .i_clk(i_clk));
Add0000000001  u_000000026B_Add0000000001(.i_data_1(matrix_r[615*12+:12]), .i_data_2(matrix_i[615*12+:12]), .o_data(c_plus_d[103][2]), .i_clk(i_clk));
Add0000000001  u_000000026C_Add0000000001(.i_data_1(matrix_r[616*12+:12]), .i_data_2(matrix_i[616*12+:12]), .o_data(c_plus_d[104][2]), .i_clk(i_clk));
Add0000000001  u_000000026D_Add0000000001(.i_data_1(matrix_r[617*12+:12]), .i_data_2(matrix_i[617*12+:12]), .o_data(c_plus_d[105][2]), .i_clk(i_clk));
Add0000000001  u_000000026E_Add0000000001(.i_data_1(matrix_r[618*12+:12]), .i_data_2(matrix_i[618*12+:12]), .o_data(c_plus_d[106][2]), .i_clk(i_clk));
Add0000000001  u_000000026F_Add0000000001(.i_data_1(matrix_r[619*12+:12]), .i_data_2(matrix_i[619*12+:12]), .o_data(c_plus_d[107][2]), .i_clk(i_clk));
Add0000000001  u_0000000270_Add0000000001(.i_data_1(matrix_r[620*12+:12]), .i_data_2(matrix_i[620*12+:12]), .o_data(c_plus_d[108][2]), .i_clk(i_clk));
Add0000000001  u_0000000271_Add0000000001(.i_data_1(matrix_r[621*12+:12]), .i_data_2(matrix_i[621*12+:12]), .o_data(c_plus_d[109][2]), .i_clk(i_clk));
Add0000000001  u_0000000272_Add0000000001(.i_data_1(matrix_r[622*12+:12]), .i_data_2(matrix_i[622*12+:12]), .o_data(c_plus_d[110][2]), .i_clk(i_clk));
Add0000000001  u_0000000273_Add0000000001(.i_data_1(matrix_r[623*12+:12]), .i_data_2(matrix_i[623*12+:12]), .o_data(c_plus_d[111][2]), .i_clk(i_clk));
Add0000000001  u_0000000274_Add0000000001(.i_data_1(matrix_r[624*12+:12]), .i_data_2(matrix_i[624*12+:12]), .o_data(c_plus_d[112][2]), .i_clk(i_clk));
Add0000000001  u_0000000275_Add0000000001(.i_data_1(matrix_r[625*12+:12]), .i_data_2(matrix_i[625*12+:12]), .o_data(c_plus_d[113][2]), .i_clk(i_clk));
Add0000000001  u_0000000276_Add0000000001(.i_data_1(matrix_r[626*12+:12]), .i_data_2(matrix_i[626*12+:12]), .o_data(c_plus_d[114][2]), .i_clk(i_clk));
Add0000000001  u_0000000277_Add0000000001(.i_data_1(matrix_r[627*12+:12]), .i_data_2(matrix_i[627*12+:12]), .o_data(c_plus_d[115][2]), .i_clk(i_clk));
Add0000000001  u_0000000278_Add0000000001(.i_data_1(matrix_r[628*12+:12]), .i_data_2(matrix_i[628*12+:12]), .o_data(c_plus_d[116][2]), .i_clk(i_clk));
Add0000000001  u_0000000279_Add0000000001(.i_data_1(matrix_r[629*12+:12]), .i_data_2(matrix_i[629*12+:12]), .o_data(c_plus_d[117][2]), .i_clk(i_clk));
Add0000000001  u_000000027A_Add0000000001(.i_data_1(matrix_r[630*12+:12]), .i_data_2(matrix_i[630*12+:12]), .o_data(c_plus_d[118][2]), .i_clk(i_clk));
Add0000000001  u_000000027B_Add0000000001(.i_data_1(matrix_r[631*12+:12]), .i_data_2(matrix_i[631*12+:12]), .o_data(c_plus_d[119][2]), .i_clk(i_clk));
Add0000000001  u_000000027C_Add0000000001(.i_data_1(matrix_r[632*12+:12]), .i_data_2(matrix_i[632*12+:12]), .o_data(c_plus_d[120][2]), .i_clk(i_clk));
Add0000000001  u_000000027D_Add0000000001(.i_data_1(matrix_r[633*12+:12]), .i_data_2(matrix_i[633*12+:12]), .o_data(c_plus_d[121][2]), .i_clk(i_clk));
Add0000000001  u_000000027E_Add0000000001(.i_data_1(matrix_r[634*12+:12]), .i_data_2(matrix_i[634*12+:12]), .o_data(c_plus_d[122][2]), .i_clk(i_clk));
Add0000000001  u_000000027F_Add0000000001(.i_data_1(matrix_r[635*12+:12]), .i_data_2(matrix_i[635*12+:12]), .o_data(c_plus_d[123][2]), .i_clk(i_clk));
Add0000000001  u_0000000280_Add0000000001(.i_data_1(matrix_r[636*12+:12]), .i_data_2(matrix_i[636*12+:12]), .o_data(c_plus_d[124][2]), .i_clk(i_clk));
Add0000000001  u_0000000281_Add0000000001(.i_data_1(matrix_r[637*12+:12]), .i_data_2(matrix_i[637*12+:12]), .o_data(c_plus_d[125][2]), .i_clk(i_clk));
Add0000000001  u_0000000282_Add0000000001(.i_data_1(matrix_r[638*12+:12]), .i_data_2(matrix_i[638*12+:12]), .o_data(c_plus_d[126][2]), .i_clk(i_clk));
Add0000000001  u_0000000283_Add0000000001(.i_data_1(matrix_r[639*12+:12]), .i_data_2(matrix_i[639*12+:12]), .o_data(c_plus_d[127][2]), .i_clk(i_clk));
Add0000000001  u_0000000284_Add0000000001(.i_data_1(matrix_r[640*12+:12]), .i_data_2(matrix_i[640*12+:12]), .o_data(c_plus_d[128][2]), .i_clk(i_clk));
Add0000000001  u_0000000285_Add0000000001(.i_data_1(matrix_r[641*12+:12]), .i_data_2(matrix_i[641*12+:12]), .o_data(c_plus_d[129][2]), .i_clk(i_clk));
Add0000000001  u_0000000286_Add0000000001(.i_data_1(matrix_r[642*12+:12]), .i_data_2(matrix_i[642*12+:12]), .o_data(c_plus_d[130][2]), .i_clk(i_clk));
Add0000000001  u_0000000287_Add0000000001(.i_data_1(matrix_r[643*12+:12]), .i_data_2(matrix_i[643*12+:12]), .o_data(c_plus_d[131][2]), .i_clk(i_clk));
Add0000000001  u_0000000288_Add0000000001(.i_data_1(matrix_r[644*12+:12]), .i_data_2(matrix_i[644*12+:12]), .o_data(c_plus_d[132][2]), .i_clk(i_clk));
Add0000000001  u_0000000289_Add0000000001(.i_data_1(matrix_r[645*12+:12]), .i_data_2(matrix_i[645*12+:12]), .o_data(c_plus_d[133][2]), .i_clk(i_clk));
Add0000000001  u_000000028A_Add0000000001(.i_data_1(matrix_r[646*12+:12]), .i_data_2(matrix_i[646*12+:12]), .o_data(c_plus_d[134][2]), .i_clk(i_clk));
Add0000000001  u_000000028B_Add0000000001(.i_data_1(matrix_r[647*12+:12]), .i_data_2(matrix_i[647*12+:12]), .o_data(c_plus_d[135][2]), .i_clk(i_clk));
Add0000000001  u_000000028C_Add0000000001(.i_data_1(matrix_r[648*12+:12]), .i_data_2(matrix_i[648*12+:12]), .o_data(c_plus_d[136][2]), .i_clk(i_clk));
Add0000000001  u_000000028D_Add0000000001(.i_data_1(matrix_r[649*12+:12]), .i_data_2(matrix_i[649*12+:12]), .o_data(c_plus_d[137][2]), .i_clk(i_clk));
Add0000000001  u_000000028E_Add0000000001(.i_data_1(matrix_r[650*12+:12]), .i_data_2(matrix_i[650*12+:12]), .o_data(c_plus_d[138][2]), .i_clk(i_clk));
Add0000000001  u_000000028F_Add0000000001(.i_data_1(matrix_r[651*12+:12]), .i_data_2(matrix_i[651*12+:12]), .o_data(c_plus_d[139][2]), .i_clk(i_clk));
Add0000000001  u_0000000290_Add0000000001(.i_data_1(matrix_r[652*12+:12]), .i_data_2(matrix_i[652*12+:12]), .o_data(c_plus_d[140][2]), .i_clk(i_clk));
Add0000000001  u_0000000291_Add0000000001(.i_data_1(matrix_r[653*12+:12]), .i_data_2(matrix_i[653*12+:12]), .o_data(c_plus_d[141][2]), .i_clk(i_clk));
Add0000000001  u_0000000292_Add0000000001(.i_data_1(matrix_r[654*12+:12]), .i_data_2(matrix_i[654*12+:12]), .o_data(c_plus_d[142][2]), .i_clk(i_clk));
Add0000000001  u_0000000293_Add0000000001(.i_data_1(matrix_r[655*12+:12]), .i_data_2(matrix_i[655*12+:12]), .o_data(c_plus_d[143][2]), .i_clk(i_clk));
Add0000000001  u_0000000294_Add0000000001(.i_data_1(matrix_r[656*12+:12]), .i_data_2(matrix_i[656*12+:12]), .o_data(c_plus_d[144][2]), .i_clk(i_clk));
Add0000000001  u_0000000295_Add0000000001(.i_data_1(matrix_r[657*12+:12]), .i_data_2(matrix_i[657*12+:12]), .o_data(c_plus_d[145][2]), .i_clk(i_clk));
Add0000000001  u_0000000296_Add0000000001(.i_data_1(matrix_r[658*12+:12]), .i_data_2(matrix_i[658*12+:12]), .o_data(c_plus_d[146][2]), .i_clk(i_clk));
Add0000000001  u_0000000297_Add0000000001(.i_data_1(matrix_r[659*12+:12]), .i_data_2(matrix_i[659*12+:12]), .o_data(c_plus_d[147][2]), .i_clk(i_clk));
Add0000000001  u_0000000298_Add0000000001(.i_data_1(matrix_r[660*12+:12]), .i_data_2(matrix_i[660*12+:12]), .o_data(c_plus_d[148][2]), .i_clk(i_clk));
Add0000000001  u_0000000299_Add0000000001(.i_data_1(matrix_r[661*12+:12]), .i_data_2(matrix_i[661*12+:12]), .o_data(c_plus_d[149][2]), .i_clk(i_clk));
Add0000000001  u_000000029A_Add0000000001(.i_data_1(matrix_r[662*12+:12]), .i_data_2(matrix_i[662*12+:12]), .o_data(c_plus_d[150][2]), .i_clk(i_clk));
Add0000000001  u_000000029B_Add0000000001(.i_data_1(matrix_r[663*12+:12]), .i_data_2(matrix_i[663*12+:12]), .o_data(c_plus_d[151][2]), .i_clk(i_clk));
Add0000000001  u_000000029C_Add0000000001(.i_data_1(matrix_r[664*12+:12]), .i_data_2(matrix_i[664*12+:12]), .o_data(c_plus_d[152][2]), .i_clk(i_clk));
Add0000000001  u_000000029D_Add0000000001(.i_data_1(matrix_r[665*12+:12]), .i_data_2(matrix_i[665*12+:12]), .o_data(c_plus_d[153][2]), .i_clk(i_clk));
Add0000000001  u_000000029E_Add0000000001(.i_data_1(matrix_r[666*12+:12]), .i_data_2(matrix_i[666*12+:12]), .o_data(c_plus_d[154][2]), .i_clk(i_clk));
Add0000000001  u_000000029F_Add0000000001(.i_data_1(matrix_r[667*12+:12]), .i_data_2(matrix_i[667*12+:12]), .o_data(c_plus_d[155][2]), .i_clk(i_clk));
Add0000000001  u_00000002A0_Add0000000001(.i_data_1(matrix_r[668*12+:12]), .i_data_2(matrix_i[668*12+:12]), .o_data(c_plus_d[156][2]), .i_clk(i_clk));
Add0000000001  u_00000002A1_Add0000000001(.i_data_1(matrix_r[669*12+:12]), .i_data_2(matrix_i[669*12+:12]), .o_data(c_plus_d[157][2]), .i_clk(i_clk));
Add0000000001  u_00000002A2_Add0000000001(.i_data_1(matrix_r[670*12+:12]), .i_data_2(matrix_i[670*12+:12]), .o_data(c_plus_d[158][2]), .i_clk(i_clk));
Add0000000001  u_00000002A3_Add0000000001(.i_data_1(matrix_r[671*12+:12]), .i_data_2(matrix_i[671*12+:12]), .o_data(c_plus_d[159][2]), .i_clk(i_clk));
Add0000000001  u_00000002A4_Add0000000001(.i_data_1(matrix_r[672*12+:12]), .i_data_2(matrix_i[672*12+:12]), .o_data(c_plus_d[160][2]), .i_clk(i_clk));
Add0000000001  u_00000002A5_Add0000000001(.i_data_1(matrix_r[673*12+:12]), .i_data_2(matrix_i[673*12+:12]), .o_data(c_plus_d[161][2]), .i_clk(i_clk));
Add0000000001  u_00000002A6_Add0000000001(.i_data_1(matrix_r[674*12+:12]), .i_data_2(matrix_i[674*12+:12]), .o_data(c_plus_d[162][2]), .i_clk(i_clk));
Add0000000001  u_00000002A7_Add0000000001(.i_data_1(matrix_r[675*12+:12]), .i_data_2(matrix_i[675*12+:12]), .o_data(c_plus_d[163][2]), .i_clk(i_clk));
Add0000000001  u_00000002A8_Add0000000001(.i_data_1(matrix_r[676*12+:12]), .i_data_2(matrix_i[676*12+:12]), .o_data(c_plus_d[164][2]), .i_clk(i_clk));
Add0000000001  u_00000002A9_Add0000000001(.i_data_1(matrix_r[677*12+:12]), .i_data_2(matrix_i[677*12+:12]), .o_data(c_plus_d[165][2]), .i_clk(i_clk));
Add0000000001  u_00000002AA_Add0000000001(.i_data_1(matrix_r[678*12+:12]), .i_data_2(matrix_i[678*12+:12]), .o_data(c_plus_d[166][2]), .i_clk(i_clk));
Add0000000001  u_00000002AB_Add0000000001(.i_data_1(matrix_r[679*12+:12]), .i_data_2(matrix_i[679*12+:12]), .o_data(c_plus_d[167][2]), .i_clk(i_clk));
Add0000000001  u_00000002AC_Add0000000001(.i_data_1(matrix_r[680*12+:12]), .i_data_2(matrix_i[680*12+:12]), .o_data(c_plus_d[168][2]), .i_clk(i_clk));
Add0000000001  u_00000002AD_Add0000000001(.i_data_1(matrix_r[681*12+:12]), .i_data_2(matrix_i[681*12+:12]), .o_data(c_plus_d[169][2]), .i_clk(i_clk));
Add0000000001  u_00000002AE_Add0000000001(.i_data_1(matrix_r[682*12+:12]), .i_data_2(matrix_i[682*12+:12]), .o_data(c_plus_d[170][2]), .i_clk(i_clk));
Add0000000001  u_00000002AF_Add0000000001(.i_data_1(matrix_r[683*12+:12]), .i_data_2(matrix_i[683*12+:12]), .o_data(c_plus_d[171][2]), .i_clk(i_clk));
Add0000000001  u_00000002B0_Add0000000001(.i_data_1(matrix_r[684*12+:12]), .i_data_2(matrix_i[684*12+:12]), .o_data(c_plus_d[172][2]), .i_clk(i_clk));
Add0000000001  u_00000002B1_Add0000000001(.i_data_1(matrix_r[685*12+:12]), .i_data_2(matrix_i[685*12+:12]), .o_data(c_plus_d[173][2]), .i_clk(i_clk));
Add0000000001  u_00000002B2_Add0000000001(.i_data_1(matrix_r[686*12+:12]), .i_data_2(matrix_i[686*12+:12]), .o_data(c_plus_d[174][2]), .i_clk(i_clk));
Add0000000001  u_00000002B3_Add0000000001(.i_data_1(matrix_r[687*12+:12]), .i_data_2(matrix_i[687*12+:12]), .o_data(c_plus_d[175][2]), .i_clk(i_clk));
Add0000000001  u_00000002B4_Add0000000001(.i_data_1(matrix_r[688*12+:12]), .i_data_2(matrix_i[688*12+:12]), .o_data(c_plus_d[176][2]), .i_clk(i_clk));
Add0000000001  u_00000002B5_Add0000000001(.i_data_1(matrix_r[689*12+:12]), .i_data_2(matrix_i[689*12+:12]), .o_data(c_plus_d[177][2]), .i_clk(i_clk));
Add0000000001  u_00000002B6_Add0000000001(.i_data_1(matrix_r[690*12+:12]), .i_data_2(matrix_i[690*12+:12]), .o_data(c_plus_d[178][2]), .i_clk(i_clk));
Add0000000001  u_00000002B7_Add0000000001(.i_data_1(matrix_r[691*12+:12]), .i_data_2(matrix_i[691*12+:12]), .o_data(c_plus_d[179][2]), .i_clk(i_clk));
Add0000000001  u_00000002B8_Add0000000001(.i_data_1(matrix_r[692*12+:12]), .i_data_2(matrix_i[692*12+:12]), .o_data(c_plus_d[180][2]), .i_clk(i_clk));
Add0000000001  u_00000002B9_Add0000000001(.i_data_1(matrix_r[693*12+:12]), .i_data_2(matrix_i[693*12+:12]), .o_data(c_plus_d[181][2]), .i_clk(i_clk));
Add0000000001  u_00000002BA_Add0000000001(.i_data_1(matrix_r[694*12+:12]), .i_data_2(matrix_i[694*12+:12]), .o_data(c_plus_d[182][2]), .i_clk(i_clk));
Add0000000001  u_00000002BB_Add0000000001(.i_data_1(matrix_r[695*12+:12]), .i_data_2(matrix_i[695*12+:12]), .o_data(c_plus_d[183][2]), .i_clk(i_clk));
Add0000000001  u_00000002BC_Add0000000001(.i_data_1(matrix_r[696*12+:12]), .i_data_2(matrix_i[696*12+:12]), .o_data(c_plus_d[184][2]), .i_clk(i_clk));
Add0000000001  u_00000002BD_Add0000000001(.i_data_1(matrix_r[697*12+:12]), .i_data_2(matrix_i[697*12+:12]), .o_data(c_plus_d[185][2]), .i_clk(i_clk));
Add0000000001  u_00000002BE_Add0000000001(.i_data_1(matrix_r[698*12+:12]), .i_data_2(matrix_i[698*12+:12]), .o_data(c_plus_d[186][2]), .i_clk(i_clk));
Add0000000001  u_00000002BF_Add0000000001(.i_data_1(matrix_r[699*12+:12]), .i_data_2(matrix_i[699*12+:12]), .o_data(c_plus_d[187][2]), .i_clk(i_clk));
Add0000000001  u_00000002C0_Add0000000001(.i_data_1(matrix_r[700*12+:12]), .i_data_2(matrix_i[700*12+:12]), .o_data(c_plus_d[188][2]), .i_clk(i_clk));
Add0000000001  u_00000002C1_Add0000000001(.i_data_1(matrix_r[701*12+:12]), .i_data_2(matrix_i[701*12+:12]), .o_data(c_plus_d[189][2]), .i_clk(i_clk));
Add0000000001  u_00000002C2_Add0000000001(.i_data_1(matrix_r[702*12+:12]), .i_data_2(matrix_i[702*12+:12]), .o_data(c_plus_d[190][2]), .i_clk(i_clk));
Add0000000001  u_00000002C3_Add0000000001(.i_data_1(matrix_r[703*12+:12]), .i_data_2(matrix_i[703*12+:12]), .o_data(c_plus_d[191][2]), .i_clk(i_clk));
Add0000000001  u_00000002C4_Add0000000001(.i_data_1(matrix_r[704*12+:12]), .i_data_2(matrix_i[704*12+:12]), .o_data(c_plus_d[192][2]), .i_clk(i_clk));
Add0000000001  u_00000002C5_Add0000000001(.i_data_1(matrix_r[705*12+:12]), .i_data_2(matrix_i[705*12+:12]), .o_data(c_plus_d[193][2]), .i_clk(i_clk));
Add0000000001  u_00000002C6_Add0000000001(.i_data_1(matrix_r[706*12+:12]), .i_data_2(matrix_i[706*12+:12]), .o_data(c_plus_d[194][2]), .i_clk(i_clk));
Add0000000001  u_00000002C7_Add0000000001(.i_data_1(matrix_r[707*12+:12]), .i_data_2(matrix_i[707*12+:12]), .o_data(c_plus_d[195][2]), .i_clk(i_clk));
Add0000000001  u_00000002C8_Add0000000001(.i_data_1(matrix_r[708*12+:12]), .i_data_2(matrix_i[708*12+:12]), .o_data(c_plus_d[196][2]), .i_clk(i_clk));
Add0000000001  u_00000002C9_Add0000000001(.i_data_1(matrix_r[709*12+:12]), .i_data_2(matrix_i[709*12+:12]), .o_data(c_plus_d[197][2]), .i_clk(i_clk));
Add0000000001  u_00000002CA_Add0000000001(.i_data_1(matrix_r[710*12+:12]), .i_data_2(matrix_i[710*12+:12]), .o_data(c_plus_d[198][2]), .i_clk(i_clk));
Add0000000001  u_00000002CB_Add0000000001(.i_data_1(matrix_r[711*12+:12]), .i_data_2(matrix_i[711*12+:12]), .o_data(c_plus_d[199][2]), .i_clk(i_clk));
Add0000000001  u_00000002CC_Add0000000001(.i_data_1(matrix_r[712*12+:12]), .i_data_2(matrix_i[712*12+:12]), .o_data(c_plus_d[200][2]), .i_clk(i_clk));
Add0000000001  u_00000002CD_Add0000000001(.i_data_1(matrix_r[713*12+:12]), .i_data_2(matrix_i[713*12+:12]), .o_data(c_plus_d[201][2]), .i_clk(i_clk));
Add0000000001  u_00000002CE_Add0000000001(.i_data_1(matrix_r[714*12+:12]), .i_data_2(matrix_i[714*12+:12]), .o_data(c_plus_d[202][2]), .i_clk(i_clk));
Add0000000001  u_00000002CF_Add0000000001(.i_data_1(matrix_r[715*12+:12]), .i_data_2(matrix_i[715*12+:12]), .o_data(c_plus_d[203][2]), .i_clk(i_clk));
Add0000000001  u_00000002D0_Add0000000001(.i_data_1(matrix_r[716*12+:12]), .i_data_2(matrix_i[716*12+:12]), .o_data(c_plus_d[204][2]), .i_clk(i_clk));
Add0000000001  u_00000002D1_Add0000000001(.i_data_1(matrix_r[717*12+:12]), .i_data_2(matrix_i[717*12+:12]), .o_data(c_plus_d[205][2]), .i_clk(i_clk));
Add0000000001  u_00000002D2_Add0000000001(.i_data_1(matrix_r[718*12+:12]), .i_data_2(matrix_i[718*12+:12]), .o_data(c_plus_d[206][2]), .i_clk(i_clk));
Add0000000001  u_00000002D3_Add0000000001(.i_data_1(matrix_r[719*12+:12]), .i_data_2(matrix_i[719*12+:12]), .o_data(c_plus_d[207][2]), .i_clk(i_clk));
Add0000000001  u_00000002D4_Add0000000001(.i_data_1(matrix_r[720*12+:12]), .i_data_2(matrix_i[720*12+:12]), .o_data(c_plus_d[208][2]), .i_clk(i_clk));
Add0000000001  u_00000002D5_Add0000000001(.i_data_1(matrix_r[721*12+:12]), .i_data_2(matrix_i[721*12+:12]), .o_data(c_plus_d[209][2]), .i_clk(i_clk));
Add0000000001  u_00000002D6_Add0000000001(.i_data_1(matrix_r[722*12+:12]), .i_data_2(matrix_i[722*12+:12]), .o_data(c_plus_d[210][2]), .i_clk(i_clk));
Add0000000001  u_00000002D7_Add0000000001(.i_data_1(matrix_r[723*12+:12]), .i_data_2(matrix_i[723*12+:12]), .o_data(c_plus_d[211][2]), .i_clk(i_clk));
Add0000000001  u_00000002D8_Add0000000001(.i_data_1(matrix_r[724*12+:12]), .i_data_2(matrix_i[724*12+:12]), .o_data(c_plus_d[212][2]), .i_clk(i_clk));
Add0000000001  u_00000002D9_Add0000000001(.i_data_1(matrix_r[725*12+:12]), .i_data_2(matrix_i[725*12+:12]), .o_data(c_plus_d[213][2]), .i_clk(i_clk));
Add0000000001  u_00000002DA_Add0000000001(.i_data_1(matrix_r[726*12+:12]), .i_data_2(matrix_i[726*12+:12]), .o_data(c_plus_d[214][2]), .i_clk(i_clk));
Add0000000001  u_00000002DB_Add0000000001(.i_data_1(matrix_r[727*12+:12]), .i_data_2(matrix_i[727*12+:12]), .o_data(c_plus_d[215][2]), .i_clk(i_clk));
Add0000000001  u_00000002DC_Add0000000001(.i_data_1(matrix_r[728*12+:12]), .i_data_2(matrix_i[728*12+:12]), .o_data(c_plus_d[216][2]), .i_clk(i_clk));
Add0000000001  u_00000002DD_Add0000000001(.i_data_1(matrix_r[729*12+:12]), .i_data_2(matrix_i[729*12+:12]), .o_data(c_plus_d[217][2]), .i_clk(i_clk));
Add0000000001  u_00000002DE_Add0000000001(.i_data_1(matrix_r[730*12+:12]), .i_data_2(matrix_i[730*12+:12]), .o_data(c_plus_d[218][2]), .i_clk(i_clk));
Add0000000001  u_00000002DF_Add0000000001(.i_data_1(matrix_r[731*12+:12]), .i_data_2(matrix_i[731*12+:12]), .o_data(c_plus_d[219][2]), .i_clk(i_clk));
Add0000000001  u_00000002E0_Add0000000001(.i_data_1(matrix_r[732*12+:12]), .i_data_2(matrix_i[732*12+:12]), .o_data(c_plus_d[220][2]), .i_clk(i_clk));
Add0000000001  u_00000002E1_Add0000000001(.i_data_1(matrix_r[733*12+:12]), .i_data_2(matrix_i[733*12+:12]), .o_data(c_plus_d[221][2]), .i_clk(i_clk));
Add0000000001  u_00000002E2_Add0000000001(.i_data_1(matrix_r[734*12+:12]), .i_data_2(matrix_i[734*12+:12]), .o_data(c_plus_d[222][2]), .i_clk(i_clk));
Add0000000001  u_00000002E3_Add0000000001(.i_data_1(matrix_r[735*12+:12]), .i_data_2(matrix_i[735*12+:12]), .o_data(c_plus_d[223][2]), .i_clk(i_clk));
Add0000000001  u_00000002E4_Add0000000001(.i_data_1(matrix_r[736*12+:12]), .i_data_2(matrix_i[736*12+:12]), .o_data(c_plus_d[224][2]), .i_clk(i_clk));
Add0000000001  u_00000002E5_Add0000000001(.i_data_1(matrix_r[737*12+:12]), .i_data_2(matrix_i[737*12+:12]), .o_data(c_plus_d[225][2]), .i_clk(i_clk));
Add0000000001  u_00000002E6_Add0000000001(.i_data_1(matrix_r[738*12+:12]), .i_data_2(matrix_i[738*12+:12]), .o_data(c_plus_d[226][2]), .i_clk(i_clk));
Add0000000001  u_00000002E7_Add0000000001(.i_data_1(matrix_r[739*12+:12]), .i_data_2(matrix_i[739*12+:12]), .o_data(c_plus_d[227][2]), .i_clk(i_clk));
Add0000000001  u_00000002E8_Add0000000001(.i_data_1(matrix_r[740*12+:12]), .i_data_2(matrix_i[740*12+:12]), .o_data(c_plus_d[228][2]), .i_clk(i_clk));
Add0000000001  u_00000002E9_Add0000000001(.i_data_1(matrix_r[741*12+:12]), .i_data_2(matrix_i[741*12+:12]), .o_data(c_plus_d[229][2]), .i_clk(i_clk));
Add0000000001  u_00000002EA_Add0000000001(.i_data_1(matrix_r[742*12+:12]), .i_data_2(matrix_i[742*12+:12]), .o_data(c_plus_d[230][2]), .i_clk(i_clk));
Add0000000001  u_00000002EB_Add0000000001(.i_data_1(matrix_r[743*12+:12]), .i_data_2(matrix_i[743*12+:12]), .o_data(c_plus_d[231][2]), .i_clk(i_clk));
Add0000000001  u_00000002EC_Add0000000001(.i_data_1(matrix_r[744*12+:12]), .i_data_2(matrix_i[744*12+:12]), .o_data(c_plus_d[232][2]), .i_clk(i_clk));
Add0000000001  u_00000002ED_Add0000000001(.i_data_1(matrix_r[745*12+:12]), .i_data_2(matrix_i[745*12+:12]), .o_data(c_plus_d[233][2]), .i_clk(i_clk));
Add0000000001  u_00000002EE_Add0000000001(.i_data_1(matrix_r[746*12+:12]), .i_data_2(matrix_i[746*12+:12]), .o_data(c_plus_d[234][2]), .i_clk(i_clk));
Add0000000001  u_00000002EF_Add0000000001(.i_data_1(matrix_r[747*12+:12]), .i_data_2(matrix_i[747*12+:12]), .o_data(c_plus_d[235][2]), .i_clk(i_clk));
Add0000000001  u_00000002F0_Add0000000001(.i_data_1(matrix_r[748*12+:12]), .i_data_2(matrix_i[748*12+:12]), .o_data(c_plus_d[236][2]), .i_clk(i_clk));
Add0000000001  u_00000002F1_Add0000000001(.i_data_1(matrix_r[749*12+:12]), .i_data_2(matrix_i[749*12+:12]), .o_data(c_plus_d[237][2]), .i_clk(i_clk));
Add0000000001  u_00000002F2_Add0000000001(.i_data_1(matrix_r[750*12+:12]), .i_data_2(matrix_i[750*12+:12]), .o_data(c_plus_d[238][2]), .i_clk(i_clk));
Add0000000001  u_00000002F3_Add0000000001(.i_data_1(matrix_r[751*12+:12]), .i_data_2(matrix_i[751*12+:12]), .o_data(c_plus_d[239][2]), .i_clk(i_clk));
Add0000000001  u_00000002F4_Add0000000001(.i_data_1(matrix_r[752*12+:12]), .i_data_2(matrix_i[752*12+:12]), .o_data(c_plus_d[240][2]), .i_clk(i_clk));
Add0000000001  u_00000002F5_Add0000000001(.i_data_1(matrix_r[753*12+:12]), .i_data_2(matrix_i[753*12+:12]), .o_data(c_plus_d[241][2]), .i_clk(i_clk));
Add0000000001  u_00000002F6_Add0000000001(.i_data_1(matrix_r[754*12+:12]), .i_data_2(matrix_i[754*12+:12]), .o_data(c_plus_d[242][2]), .i_clk(i_clk));
Add0000000001  u_00000002F7_Add0000000001(.i_data_1(matrix_r[755*12+:12]), .i_data_2(matrix_i[755*12+:12]), .o_data(c_plus_d[243][2]), .i_clk(i_clk));
Add0000000001  u_00000002F8_Add0000000001(.i_data_1(matrix_r[756*12+:12]), .i_data_2(matrix_i[756*12+:12]), .o_data(c_plus_d[244][2]), .i_clk(i_clk));
Add0000000001  u_00000002F9_Add0000000001(.i_data_1(matrix_r[757*12+:12]), .i_data_2(matrix_i[757*12+:12]), .o_data(c_plus_d[245][2]), .i_clk(i_clk));
Add0000000001  u_00000002FA_Add0000000001(.i_data_1(matrix_r[758*12+:12]), .i_data_2(matrix_i[758*12+:12]), .o_data(c_plus_d[246][2]), .i_clk(i_clk));
Add0000000001  u_00000002FB_Add0000000001(.i_data_1(matrix_r[759*12+:12]), .i_data_2(matrix_i[759*12+:12]), .o_data(c_plus_d[247][2]), .i_clk(i_clk));
Add0000000001  u_00000002FC_Add0000000001(.i_data_1(matrix_r[760*12+:12]), .i_data_2(matrix_i[760*12+:12]), .o_data(c_plus_d[248][2]), .i_clk(i_clk));
Add0000000001  u_00000002FD_Add0000000001(.i_data_1(matrix_r[761*12+:12]), .i_data_2(matrix_i[761*12+:12]), .o_data(c_plus_d[249][2]), .i_clk(i_clk));
Add0000000001  u_00000002FE_Add0000000001(.i_data_1(matrix_r[762*12+:12]), .i_data_2(matrix_i[762*12+:12]), .o_data(c_plus_d[250][2]), .i_clk(i_clk));
Add0000000001  u_00000002FF_Add0000000001(.i_data_1(matrix_r[763*12+:12]), .i_data_2(matrix_i[763*12+:12]), .o_data(c_plus_d[251][2]), .i_clk(i_clk));
Add0000000001  u_0000000300_Add0000000001(.i_data_1(matrix_r[764*12+:12]), .i_data_2(matrix_i[764*12+:12]), .o_data(c_plus_d[252][2]), .i_clk(i_clk));
Add0000000001  u_0000000301_Add0000000001(.i_data_1(matrix_r[765*12+:12]), .i_data_2(matrix_i[765*12+:12]), .o_data(c_plus_d[253][2]), .i_clk(i_clk));
Add0000000001  u_0000000302_Add0000000001(.i_data_1(matrix_r[766*12+:12]), .i_data_2(matrix_i[766*12+:12]), .o_data(c_plus_d[254][2]), .i_clk(i_clk));
Add0000000001  u_0000000303_Add0000000001(.i_data_1(matrix_r[767*12+:12]), .i_data_2(matrix_i[767*12+:12]), .o_data(c_plus_d[255][2]), .i_clk(i_clk));
Add0000000001  u_0000000304_Add0000000001(.i_data_1(vector_r[3*12+:12]), .i_data_2(vector_i[3*12+:12]), .o_data(a_plus_b[3]), .i_clk(i_clk));
Sub0000000001  u_0000000004_Sub0000000001(.i_data_1(vector_i[3*12+:12]), .i_data_2(vector_r[3*12+:12]), .o_data(b_minus_a[3]), .i_clk(i_clk));
Add0000000001  u_0000000305_Add0000000001(.i_data_1(matrix_r[768*12+:12]), .i_data_2(matrix_i[768*12+:12]), .o_data(c_plus_d[0][3]), .i_clk(i_clk));
Add0000000001  u_0000000306_Add0000000001(.i_data_1(matrix_r[769*12+:12]), .i_data_2(matrix_i[769*12+:12]), .o_data(c_plus_d[1][3]), .i_clk(i_clk));
Add0000000001  u_0000000307_Add0000000001(.i_data_1(matrix_r[770*12+:12]), .i_data_2(matrix_i[770*12+:12]), .o_data(c_plus_d[2][3]), .i_clk(i_clk));
Add0000000001  u_0000000308_Add0000000001(.i_data_1(matrix_r[771*12+:12]), .i_data_2(matrix_i[771*12+:12]), .o_data(c_plus_d[3][3]), .i_clk(i_clk));
Add0000000001  u_0000000309_Add0000000001(.i_data_1(matrix_r[772*12+:12]), .i_data_2(matrix_i[772*12+:12]), .o_data(c_plus_d[4][3]), .i_clk(i_clk));
Add0000000001  u_000000030A_Add0000000001(.i_data_1(matrix_r[773*12+:12]), .i_data_2(matrix_i[773*12+:12]), .o_data(c_plus_d[5][3]), .i_clk(i_clk));
Add0000000001  u_000000030B_Add0000000001(.i_data_1(matrix_r[774*12+:12]), .i_data_2(matrix_i[774*12+:12]), .o_data(c_plus_d[6][3]), .i_clk(i_clk));
Add0000000001  u_000000030C_Add0000000001(.i_data_1(matrix_r[775*12+:12]), .i_data_2(matrix_i[775*12+:12]), .o_data(c_plus_d[7][3]), .i_clk(i_clk));
Add0000000001  u_000000030D_Add0000000001(.i_data_1(matrix_r[776*12+:12]), .i_data_2(matrix_i[776*12+:12]), .o_data(c_plus_d[8][3]), .i_clk(i_clk));
Add0000000001  u_000000030E_Add0000000001(.i_data_1(matrix_r[777*12+:12]), .i_data_2(matrix_i[777*12+:12]), .o_data(c_plus_d[9][3]), .i_clk(i_clk));
Add0000000001  u_000000030F_Add0000000001(.i_data_1(matrix_r[778*12+:12]), .i_data_2(matrix_i[778*12+:12]), .o_data(c_plus_d[10][3]), .i_clk(i_clk));
Add0000000001  u_0000000310_Add0000000001(.i_data_1(matrix_r[779*12+:12]), .i_data_2(matrix_i[779*12+:12]), .o_data(c_plus_d[11][3]), .i_clk(i_clk));
Add0000000001  u_0000000311_Add0000000001(.i_data_1(matrix_r[780*12+:12]), .i_data_2(matrix_i[780*12+:12]), .o_data(c_plus_d[12][3]), .i_clk(i_clk));
Add0000000001  u_0000000312_Add0000000001(.i_data_1(matrix_r[781*12+:12]), .i_data_2(matrix_i[781*12+:12]), .o_data(c_plus_d[13][3]), .i_clk(i_clk));
Add0000000001  u_0000000313_Add0000000001(.i_data_1(matrix_r[782*12+:12]), .i_data_2(matrix_i[782*12+:12]), .o_data(c_plus_d[14][3]), .i_clk(i_clk));
Add0000000001  u_0000000314_Add0000000001(.i_data_1(matrix_r[783*12+:12]), .i_data_2(matrix_i[783*12+:12]), .o_data(c_plus_d[15][3]), .i_clk(i_clk));
Add0000000001  u_0000000315_Add0000000001(.i_data_1(matrix_r[784*12+:12]), .i_data_2(matrix_i[784*12+:12]), .o_data(c_plus_d[16][3]), .i_clk(i_clk));
Add0000000001  u_0000000316_Add0000000001(.i_data_1(matrix_r[785*12+:12]), .i_data_2(matrix_i[785*12+:12]), .o_data(c_plus_d[17][3]), .i_clk(i_clk));
Add0000000001  u_0000000317_Add0000000001(.i_data_1(matrix_r[786*12+:12]), .i_data_2(matrix_i[786*12+:12]), .o_data(c_plus_d[18][3]), .i_clk(i_clk));
Add0000000001  u_0000000318_Add0000000001(.i_data_1(matrix_r[787*12+:12]), .i_data_2(matrix_i[787*12+:12]), .o_data(c_plus_d[19][3]), .i_clk(i_clk));
Add0000000001  u_0000000319_Add0000000001(.i_data_1(matrix_r[788*12+:12]), .i_data_2(matrix_i[788*12+:12]), .o_data(c_plus_d[20][3]), .i_clk(i_clk));
Add0000000001  u_000000031A_Add0000000001(.i_data_1(matrix_r[789*12+:12]), .i_data_2(matrix_i[789*12+:12]), .o_data(c_plus_d[21][3]), .i_clk(i_clk));
Add0000000001  u_000000031B_Add0000000001(.i_data_1(matrix_r[790*12+:12]), .i_data_2(matrix_i[790*12+:12]), .o_data(c_plus_d[22][3]), .i_clk(i_clk));
Add0000000001  u_000000031C_Add0000000001(.i_data_1(matrix_r[791*12+:12]), .i_data_2(matrix_i[791*12+:12]), .o_data(c_plus_d[23][3]), .i_clk(i_clk));
Add0000000001  u_000000031D_Add0000000001(.i_data_1(matrix_r[792*12+:12]), .i_data_2(matrix_i[792*12+:12]), .o_data(c_plus_d[24][3]), .i_clk(i_clk));
Add0000000001  u_000000031E_Add0000000001(.i_data_1(matrix_r[793*12+:12]), .i_data_2(matrix_i[793*12+:12]), .o_data(c_plus_d[25][3]), .i_clk(i_clk));
Add0000000001  u_000000031F_Add0000000001(.i_data_1(matrix_r[794*12+:12]), .i_data_2(matrix_i[794*12+:12]), .o_data(c_plus_d[26][3]), .i_clk(i_clk));
Add0000000001  u_0000000320_Add0000000001(.i_data_1(matrix_r[795*12+:12]), .i_data_2(matrix_i[795*12+:12]), .o_data(c_plus_d[27][3]), .i_clk(i_clk));
Add0000000001  u_0000000321_Add0000000001(.i_data_1(matrix_r[796*12+:12]), .i_data_2(matrix_i[796*12+:12]), .o_data(c_plus_d[28][3]), .i_clk(i_clk));
Add0000000001  u_0000000322_Add0000000001(.i_data_1(matrix_r[797*12+:12]), .i_data_2(matrix_i[797*12+:12]), .o_data(c_plus_d[29][3]), .i_clk(i_clk));
Add0000000001  u_0000000323_Add0000000001(.i_data_1(matrix_r[798*12+:12]), .i_data_2(matrix_i[798*12+:12]), .o_data(c_plus_d[30][3]), .i_clk(i_clk));
Add0000000001  u_0000000324_Add0000000001(.i_data_1(matrix_r[799*12+:12]), .i_data_2(matrix_i[799*12+:12]), .o_data(c_plus_d[31][3]), .i_clk(i_clk));
Add0000000001  u_0000000325_Add0000000001(.i_data_1(matrix_r[800*12+:12]), .i_data_2(matrix_i[800*12+:12]), .o_data(c_plus_d[32][3]), .i_clk(i_clk));
Add0000000001  u_0000000326_Add0000000001(.i_data_1(matrix_r[801*12+:12]), .i_data_2(matrix_i[801*12+:12]), .o_data(c_plus_d[33][3]), .i_clk(i_clk));
Add0000000001  u_0000000327_Add0000000001(.i_data_1(matrix_r[802*12+:12]), .i_data_2(matrix_i[802*12+:12]), .o_data(c_plus_d[34][3]), .i_clk(i_clk));
Add0000000001  u_0000000328_Add0000000001(.i_data_1(matrix_r[803*12+:12]), .i_data_2(matrix_i[803*12+:12]), .o_data(c_plus_d[35][3]), .i_clk(i_clk));
Add0000000001  u_0000000329_Add0000000001(.i_data_1(matrix_r[804*12+:12]), .i_data_2(matrix_i[804*12+:12]), .o_data(c_plus_d[36][3]), .i_clk(i_clk));
Add0000000001  u_000000032A_Add0000000001(.i_data_1(matrix_r[805*12+:12]), .i_data_2(matrix_i[805*12+:12]), .o_data(c_plus_d[37][3]), .i_clk(i_clk));
Add0000000001  u_000000032B_Add0000000001(.i_data_1(matrix_r[806*12+:12]), .i_data_2(matrix_i[806*12+:12]), .o_data(c_plus_d[38][3]), .i_clk(i_clk));
Add0000000001  u_000000032C_Add0000000001(.i_data_1(matrix_r[807*12+:12]), .i_data_2(matrix_i[807*12+:12]), .o_data(c_plus_d[39][3]), .i_clk(i_clk));
Add0000000001  u_000000032D_Add0000000001(.i_data_1(matrix_r[808*12+:12]), .i_data_2(matrix_i[808*12+:12]), .o_data(c_plus_d[40][3]), .i_clk(i_clk));
Add0000000001  u_000000032E_Add0000000001(.i_data_1(matrix_r[809*12+:12]), .i_data_2(matrix_i[809*12+:12]), .o_data(c_plus_d[41][3]), .i_clk(i_clk));
Add0000000001  u_000000032F_Add0000000001(.i_data_1(matrix_r[810*12+:12]), .i_data_2(matrix_i[810*12+:12]), .o_data(c_plus_d[42][3]), .i_clk(i_clk));
Add0000000001  u_0000000330_Add0000000001(.i_data_1(matrix_r[811*12+:12]), .i_data_2(matrix_i[811*12+:12]), .o_data(c_plus_d[43][3]), .i_clk(i_clk));
Add0000000001  u_0000000331_Add0000000001(.i_data_1(matrix_r[812*12+:12]), .i_data_2(matrix_i[812*12+:12]), .o_data(c_plus_d[44][3]), .i_clk(i_clk));
Add0000000001  u_0000000332_Add0000000001(.i_data_1(matrix_r[813*12+:12]), .i_data_2(matrix_i[813*12+:12]), .o_data(c_plus_d[45][3]), .i_clk(i_clk));
Add0000000001  u_0000000333_Add0000000001(.i_data_1(matrix_r[814*12+:12]), .i_data_2(matrix_i[814*12+:12]), .o_data(c_plus_d[46][3]), .i_clk(i_clk));
Add0000000001  u_0000000334_Add0000000001(.i_data_1(matrix_r[815*12+:12]), .i_data_2(matrix_i[815*12+:12]), .o_data(c_plus_d[47][3]), .i_clk(i_clk));
Add0000000001  u_0000000335_Add0000000001(.i_data_1(matrix_r[816*12+:12]), .i_data_2(matrix_i[816*12+:12]), .o_data(c_plus_d[48][3]), .i_clk(i_clk));
Add0000000001  u_0000000336_Add0000000001(.i_data_1(matrix_r[817*12+:12]), .i_data_2(matrix_i[817*12+:12]), .o_data(c_plus_d[49][3]), .i_clk(i_clk));
Add0000000001  u_0000000337_Add0000000001(.i_data_1(matrix_r[818*12+:12]), .i_data_2(matrix_i[818*12+:12]), .o_data(c_plus_d[50][3]), .i_clk(i_clk));
Add0000000001  u_0000000338_Add0000000001(.i_data_1(matrix_r[819*12+:12]), .i_data_2(matrix_i[819*12+:12]), .o_data(c_plus_d[51][3]), .i_clk(i_clk));
Add0000000001  u_0000000339_Add0000000001(.i_data_1(matrix_r[820*12+:12]), .i_data_2(matrix_i[820*12+:12]), .o_data(c_plus_d[52][3]), .i_clk(i_clk));
Add0000000001  u_000000033A_Add0000000001(.i_data_1(matrix_r[821*12+:12]), .i_data_2(matrix_i[821*12+:12]), .o_data(c_plus_d[53][3]), .i_clk(i_clk));
Add0000000001  u_000000033B_Add0000000001(.i_data_1(matrix_r[822*12+:12]), .i_data_2(matrix_i[822*12+:12]), .o_data(c_plus_d[54][3]), .i_clk(i_clk));
Add0000000001  u_000000033C_Add0000000001(.i_data_1(matrix_r[823*12+:12]), .i_data_2(matrix_i[823*12+:12]), .o_data(c_plus_d[55][3]), .i_clk(i_clk));
Add0000000001  u_000000033D_Add0000000001(.i_data_1(matrix_r[824*12+:12]), .i_data_2(matrix_i[824*12+:12]), .o_data(c_plus_d[56][3]), .i_clk(i_clk));
Add0000000001  u_000000033E_Add0000000001(.i_data_1(matrix_r[825*12+:12]), .i_data_2(matrix_i[825*12+:12]), .o_data(c_plus_d[57][3]), .i_clk(i_clk));
Add0000000001  u_000000033F_Add0000000001(.i_data_1(matrix_r[826*12+:12]), .i_data_2(matrix_i[826*12+:12]), .o_data(c_plus_d[58][3]), .i_clk(i_clk));
Add0000000001  u_0000000340_Add0000000001(.i_data_1(matrix_r[827*12+:12]), .i_data_2(matrix_i[827*12+:12]), .o_data(c_plus_d[59][3]), .i_clk(i_clk));
Add0000000001  u_0000000341_Add0000000001(.i_data_1(matrix_r[828*12+:12]), .i_data_2(matrix_i[828*12+:12]), .o_data(c_plus_d[60][3]), .i_clk(i_clk));
Add0000000001  u_0000000342_Add0000000001(.i_data_1(matrix_r[829*12+:12]), .i_data_2(matrix_i[829*12+:12]), .o_data(c_plus_d[61][3]), .i_clk(i_clk));
Add0000000001  u_0000000343_Add0000000001(.i_data_1(matrix_r[830*12+:12]), .i_data_2(matrix_i[830*12+:12]), .o_data(c_plus_d[62][3]), .i_clk(i_clk));
Add0000000001  u_0000000344_Add0000000001(.i_data_1(matrix_r[831*12+:12]), .i_data_2(matrix_i[831*12+:12]), .o_data(c_plus_d[63][3]), .i_clk(i_clk));
Add0000000001  u_0000000345_Add0000000001(.i_data_1(matrix_r[832*12+:12]), .i_data_2(matrix_i[832*12+:12]), .o_data(c_plus_d[64][3]), .i_clk(i_clk));
Add0000000001  u_0000000346_Add0000000001(.i_data_1(matrix_r[833*12+:12]), .i_data_2(matrix_i[833*12+:12]), .o_data(c_plus_d[65][3]), .i_clk(i_clk));
Add0000000001  u_0000000347_Add0000000001(.i_data_1(matrix_r[834*12+:12]), .i_data_2(matrix_i[834*12+:12]), .o_data(c_plus_d[66][3]), .i_clk(i_clk));
Add0000000001  u_0000000348_Add0000000001(.i_data_1(matrix_r[835*12+:12]), .i_data_2(matrix_i[835*12+:12]), .o_data(c_plus_d[67][3]), .i_clk(i_clk));
Add0000000001  u_0000000349_Add0000000001(.i_data_1(matrix_r[836*12+:12]), .i_data_2(matrix_i[836*12+:12]), .o_data(c_plus_d[68][3]), .i_clk(i_clk));
Add0000000001  u_000000034A_Add0000000001(.i_data_1(matrix_r[837*12+:12]), .i_data_2(matrix_i[837*12+:12]), .o_data(c_plus_d[69][3]), .i_clk(i_clk));
Add0000000001  u_000000034B_Add0000000001(.i_data_1(matrix_r[838*12+:12]), .i_data_2(matrix_i[838*12+:12]), .o_data(c_plus_d[70][3]), .i_clk(i_clk));
Add0000000001  u_000000034C_Add0000000001(.i_data_1(matrix_r[839*12+:12]), .i_data_2(matrix_i[839*12+:12]), .o_data(c_plus_d[71][3]), .i_clk(i_clk));
Add0000000001  u_000000034D_Add0000000001(.i_data_1(matrix_r[840*12+:12]), .i_data_2(matrix_i[840*12+:12]), .o_data(c_plus_d[72][3]), .i_clk(i_clk));
Add0000000001  u_000000034E_Add0000000001(.i_data_1(matrix_r[841*12+:12]), .i_data_2(matrix_i[841*12+:12]), .o_data(c_plus_d[73][3]), .i_clk(i_clk));
Add0000000001  u_000000034F_Add0000000001(.i_data_1(matrix_r[842*12+:12]), .i_data_2(matrix_i[842*12+:12]), .o_data(c_plus_d[74][3]), .i_clk(i_clk));
Add0000000001  u_0000000350_Add0000000001(.i_data_1(matrix_r[843*12+:12]), .i_data_2(matrix_i[843*12+:12]), .o_data(c_plus_d[75][3]), .i_clk(i_clk));
Add0000000001  u_0000000351_Add0000000001(.i_data_1(matrix_r[844*12+:12]), .i_data_2(matrix_i[844*12+:12]), .o_data(c_plus_d[76][3]), .i_clk(i_clk));
Add0000000001  u_0000000352_Add0000000001(.i_data_1(matrix_r[845*12+:12]), .i_data_2(matrix_i[845*12+:12]), .o_data(c_plus_d[77][3]), .i_clk(i_clk));
Add0000000001  u_0000000353_Add0000000001(.i_data_1(matrix_r[846*12+:12]), .i_data_2(matrix_i[846*12+:12]), .o_data(c_plus_d[78][3]), .i_clk(i_clk));
Add0000000001  u_0000000354_Add0000000001(.i_data_1(matrix_r[847*12+:12]), .i_data_2(matrix_i[847*12+:12]), .o_data(c_plus_d[79][3]), .i_clk(i_clk));
Add0000000001  u_0000000355_Add0000000001(.i_data_1(matrix_r[848*12+:12]), .i_data_2(matrix_i[848*12+:12]), .o_data(c_plus_d[80][3]), .i_clk(i_clk));
Add0000000001  u_0000000356_Add0000000001(.i_data_1(matrix_r[849*12+:12]), .i_data_2(matrix_i[849*12+:12]), .o_data(c_plus_d[81][3]), .i_clk(i_clk));
Add0000000001  u_0000000357_Add0000000001(.i_data_1(matrix_r[850*12+:12]), .i_data_2(matrix_i[850*12+:12]), .o_data(c_plus_d[82][3]), .i_clk(i_clk));
Add0000000001  u_0000000358_Add0000000001(.i_data_1(matrix_r[851*12+:12]), .i_data_2(matrix_i[851*12+:12]), .o_data(c_plus_d[83][3]), .i_clk(i_clk));
Add0000000001  u_0000000359_Add0000000001(.i_data_1(matrix_r[852*12+:12]), .i_data_2(matrix_i[852*12+:12]), .o_data(c_plus_d[84][3]), .i_clk(i_clk));
Add0000000001  u_000000035A_Add0000000001(.i_data_1(matrix_r[853*12+:12]), .i_data_2(matrix_i[853*12+:12]), .o_data(c_plus_d[85][3]), .i_clk(i_clk));
Add0000000001  u_000000035B_Add0000000001(.i_data_1(matrix_r[854*12+:12]), .i_data_2(matrix_i[854*12+:12]), .o_data(c_plus_d[86][3]), .i_clk(i_clk));
Add0000000001  u_000000035C_Add0000000001(.i_data_1(matrix_r[855*12+:12]), .i_data_2(matrix_i[855*12+:12]), .o_data(c_plus_d[87][3]), .i_clk(i_clk));
Add0000000001  u_000000035D_Add0000000001(.i_data_1(matrix_r[856*12+:12]), .i_data_2(matrix_i[856*12+:12]), .o_data(c_plus_d[88][3]), .i_clk(i_clk));
Add0000000001  u_000000035E_Add0000000001(.i_data_1(matrix_r[857*12+:12]), .i_data_2(matrix_i[857*12+:12]), .o_data(c_plus_d[89][3]), .i_clk(i_clk));
Add0000000001  u_000000035F_Add0000000001(.i_data_1(matrix_r[858*12+:12]), .i_data_2(matrix_i[858*12+:12]), .o_data(c_plus_d[90][3]), .i_clk(i_clk));
Add0000000001  u_0000000360_Add0000000001(.i_data_1(matrix_r[859*12+:12]), .i_data_2(matrix_i[859*12+:12]), .o_data(c_plus_d[91][3]), .i_clk(i_clk));
Add0000000001  u_0000000361_Add0000000001(.i_data_1(matrix_r[860*12+:12]), .i_data_2(matrix_i[860*12+:12]), .o_data(c_plus_d[92][3]), .i_clk(i_clk));
Add0000000001  u_0000000362_Add0000000001(.i_data_1(matrix_r[861*12+:12]), .i_data_2(matrix_i[861*12+:12]), .o_data(c_plus_d[93][3]), .i_clk(i_clk));
Add0000000001  u_0000000363_Add0000000001(.i_data_1(matrix_r[862*12+:12]), .i_data_2(matrix_i[862*12+:12]), .o_data(c_plus_d[94][3]), .i_clk(i_clk));
Add0000000001  u_0000000364_Add0000000001(.i_data_1(matrix_r[863*12+:12]), .i_data_2(matrix_i[863*12+:12]), .o_data(c_plus_d[95][3]), .i_clk(i_clk));
Add0000000001  u_0000000365_Add0000000001(.i_data_1(matrix_r[864*12+:12]), .i_data_2(matrix_i[864*12+:12]), .o_data(c_plus_d[96][3]), .i_clk(i_clk));
Add0000000001  u_0000000366_Add0000000001(.i_data_1(matrix_r[865*12+:12]), .i_data_2(matrix_i[865*12+:12]), .o_data(c_plus_d[97][3]), .i_clk(i_clk));
Add0000000001  u_0000000367_Add0000000001(.i_data_1(matrix_r[866*12+:12]), .i_data_2(matrix_i[866*12+:12]), .o_data(c_plus_d[98][3]), .i_clk(i_clk));
Add0000000001  u_0000000368_Add0000000001(.i_data_1(matrix_r[867*12+:12]), .i_data_2(matrix_i[867*12+:12]), .o_data(c_plus_d[99][3]), .i_clk(i_clk));
Add0000000001  u_0000000369_Add0000000001(.i_data_1(matrix_r[868*12+:12]), .i_data_2(matrix_i[868*12+:12]), .o_data(c_plus_d[100][3]), .i_clk(i_clk));
Add0000000001  u_000000036A_Add0000000001(.i_data_1(matrix_r[869*12+:12]), .i_data_2(matrix_i[869*12+:12]), .o_data(c_plus_d[101][3]), .i_clk(i_clk));
Add0000000001  u_000000036B_Add0000000001(.i_data_1(matrix_r[870*12+:12]), .i_data_2(matrix_i[870*12+:12]), .o_data(c_plus_d[102][3]), .i_clk(i_clk));
Add0000000001  u_000000036C_Add0000000001(.i_data_1(matrix_r[871*12+:12]), .i_data_2(matrix_i[871*12+:12]), .o_data(c_plus_d[103][3]), .i_clk(i_clk));
Add0000000001  u_000000036D_Add0000000001(.i_data_1(matrix_r[872*12+:12]), .i_data_2(matrix_i[872*12+:12]), .o_data(c_plus_d[104][3]), .i_clk(i_clk));
Add0000000001  u_000000036E_Add0000000001(.i_data_1(matrix_r[873*12+:12]), .i_data_2(matrix_i[873*12+:12]), .o_data(c_plus_d[105][3]), .i_clk(i_clk));
Add0000000001  u_000000036F_Add0000000001(.i_data_1(matrix_r[874*12+:12]), .i_data_2(matrix_i[874*12+:12]), .o_data(c_plus_d[106][3]), .i_clk(i_clk));
Add0000000001  u_0000000370_Add0000000001(.i_data_1(matrix_r[875*12+:12]), .i_data_2(matrix_i[875*12+:12]), .o_data(c_plus_d[107][3]), .i_clk(i_clk));
Add0000000001  u_0000000371_Add0000000001(.i_data_1(matrix_r[876*12+:12]), .i_data_2(matrix_i[876*12+:12]), .o_data(c_plus_d[108][3]), .i_clk(i_clk));
Add0000000001  u_0000000372_Add0000000001(.i_data_1(matrix_r[877*12+:12]), .i_data_2(matrix_i[877*12+:12]), .o_data(c_plus_d[109][3]), .i_clk(i_clk));
Add0000000001  u_0000000373_Add0000000001(.i_data_1(matrix_r[878*12+:12]), .i_data_2(matrix_i[878*12+:12]), .o_data(c_plus_d[110][3]), .i_clk(i_clk));
Add0000000001  u_0000000374_Add0000000001(.i_data_1(matrix_r[879*12+:12]), .i_data_2(matrix_i[879*12+:12]), .o_data(c_plus_d[111][3]), .i_clk(i_clk));
Add0000000001  u_0000000375_Add0000000001(.i_data_1(matrix_r[880*12+:12]), .i_data_2(matrix_i[880*12+:12]), .o_data(c_plus_d[112][3]), .i_clk(i_clk));
Add0000000001  u_0000000376_Add0000000001(.i_data_1(matrix_r[881*12+:12]), .i_data_2(matrix_i[881*12+:12]), .o_data(c_plus_d[113][3]), .i_clk(i_clk));
Add0000000001  u_0000000377_Add0000000001(.i_data_1(matrix_r[882*12+:12]), .i_data_2(matrix_i[882*12+:12]), .o_data(c_plus_d[114][3]), .i_clk(i_clk));
Add0000000001  u_0000000378_Add0000000001(.i_data_1(matrix_r[883*12+:12]), .i_data_2(matrix_i[883*12+:12]), .o_data(c_plus_d[115][3]), .i_clk(i_clk));
Add0000000001  u_0000000379_Add0000000001(.i_data_1(matrix_r[884*12+:12]), .i_data_2(matrix_i[884*12+:12]), .o_data(c_plus_d[116][3]), .i_clk(i_clk));
Add0000000001  u_000000037A_Add0000000001(.i_data_1(matrix_r[885*12+:12]), .i_data_2(matrix_i[885*12+:12]), .o_data(c_plus_d[117][3]), .i_clk(i_clk));
Add0000000001  u_000000037B_Add0000000001(.i_data_1(matrix_r[886*12+:12]), .i_data_2(matrix_i[886*12+:12]), .o_data(c_plus_d[118][3]), .i_clk(i_clk));
Add0000000001  u_000000037C_Add0000000001(.i_data_1(matrix_r[887*12+:12]), .i_data_2(matrix_i[887*12+:12]), .o_data(c_plus_d[119][3]), .i_clk(i_clk));
Add0000000001  u_000000037D_Add0000000001(.i_data_1(matrix_r[888*12+:12]), .i_data_2(matrix_i[888*12+:12]), .o_data(c_plus_d[120][3]), .i_clk(i_clk));
Add0000000001  u_000000037E_Add0000000001(.i_data_1(matrix_r[889*12+:12]), .i_data_2(matrix_i[889*12+:12]), .o_data(c_plus_d[121][3]), .i_clk(i_clk));
Add0000000001  u_000000037F_Add0000000001(.i_data_1(matrix_r[890*12+:12]), .i_data_2(matrix_i[890*12+:12]), .o_data(c_plus_d[122][3]), .i_clk(i_clk));
Add0000000001  u_0000000380_Add0000000001(.i_data_1(matrix_r[891*12+:12]), .i_data_2(matrix_i[891*12+:12]), .o_data(c_plus_d[123][3]), .i_clk(i_clk));
Add0000000001  u_0000000381_Add0000000001(.i_data_1(matrix_r[892*12+:12]), .i_data_2(matrix_i[892*12+:12]), .o_data(c_plus_d[124][3]), .i_clk(i_clk));
Add0000000001  u_0000000382_Add0000000001(.i_data_1(matrix_r[893*12+:12]), .i_data_2(matrix_i[893*12+:12]), .o_data(c_plus_d[125][3]), .i_clk(i_clk));
Add0000000001  u_0000000383_Add0000000001(.i_data_1(matrix_r[894*12+:12]), .i_data_2(matrix_i[894*12+:12]), .o_data(c_plus_d[126][3]), .i_clk(i_clk));
Add0000000001  u_0000000384_Add0000000001(.i_data_1(matrix_r[895*12+:12]), .i_data_2(matrix_i[895*12+:12]), .o_data(c_plus_d[127][3]), .i_clk(i_clk));
Add0000000001  u_0000000385_Add0000000001(.i_data_1(matrix_r[896*12+:12]), .i_data_2(matrix_i[896*12+:12]), .o_data(c_plus_d[128][3]), .i_clk(i_clk));
Add0000000001  u_0000000386_Add0000000001(.i_data_1(matrix_r[897*12+:12]), .i_data_2(matrix_i[897*12+:12]), .o_data(c_plus_d[129][3]), .i_clk(i_clk));
Add0000000001  u_0000000387_Add0000000001(.i_data_1(matrix_r[898*12+:12]), .i_data_2(matrix_i[898*12+:12]), .o_data(c_plus_d[130][3]), .i_clk(i_clk));
Add0000000001  u_0000000388_Add0000000001(.i_data_1(matrix_r[899*12+:12]), .i_data_2(matrix_i[899*12+:12]), .o_data(c_plus_d[131][3]), .i_clk(i_clk));
Add0000000001  u_0000000389_Add0000000001(.i_data_1(matrix_r[900*12+:12]), .i_data_2(matrix_i[900*12+:12]), .o_data(c_plus_d[132][3]), .i_clk(i_clk));
Add0000000001  u_000000038A_Add0000000001(.i_data_1(matrix_r[901*12+:12]), .i_data_2(matrix_i[901*12+:12]), .o_data(c_plus_d[133][3]), .i_clk(i_clk));
Add0000000001  u_000000038B_Add0000000001(.i_data_1(matrix_r[902*12+:12]), .i_data_2(matrix_i[902*12+:12]), .o_data(c_plus_d[134][3]), .i_clk(i_clk));
Add0000000001  u_000000038C_Add0000000001(.i_data_1(matrix_r[903*12+:12]), .i_data_2(matrix_i[903*12+:12]), .o_data(c_plus_d[135][3]), .i_clk(i_clk));
Add0000000001  u_000000038D_Add0000000001(.i_data_1(matrix_r[904*12+:12]), .i_data_2(matrix_i[904*12+:12]), .o_data(c_plus_d[136][3]), .i_clk(i_clk));
Add0000000001  u_000000038E_Add0000000001(.i_data_1(matrix_r[905*12+:12]), .i_data_2(matrix_i[905*12+:12]), .o_data(c_plus_d[137][3]), .i_clk(i_clk));
Add0000000001  u_000000038F_Add0000000001(.i_data_1(matrix_r[906*12+:12]), .i_data_2(matrix_i[906*12+:12]), .o_data(c_plus_d[138][3]), .i_clk(i_clk));
Add0000000001  u_0000000390_Add0000000001(.i_data_1(matrix_r[907*12+:12]), .i_data_2(matrix_i[907*12+:12]), .o_data(c_plus_d[139][3]), .i_clk(i_clk));
Add0000000001  u_0000000391_Add0000000001(.i_data_1(matrix_r[908*12+:12]), .i_data_2(matrix_i[908*12+:12]), .o_data(c_plus_d[140][3]), .i_clk(i_clk));
Add0000000001  u_0000000392_Add0000000001(.i_data_1(matrix_r[909*12+:12]), .i_data_2(matrix_i[909*12+:12]), .o_data(c_plus_d[141][3]), .i_clk(i_clk));
Add0000000001  u_0000000393_Add0000000001(.i_data_1(matrix_r[910*12+:12]), .i_data_2(matrix_i[910*12+:12]), .o_data(c_plus_d[142][3]), .i_clk(i_clk));
Add0000000001  u_0000000394_Add0000000001(.i_data_1(matrix_r[911*12+:12]), .i_data_2(matrix_i[911*12+:12]), .o_data(c_plus_d[143][3]), .i_clk(i_clk));
Add0000000001  u_0000000395_Add0000000001(.i_data_1(matrix_r[912*12+:12]), .i_data_2(matrix_i[912*12+:12]), .o_data(c_plus_d[144][3]), .i_clk(i_clk));
Add0000000001  u_0000000396_Add0000000001(.i_data_1(matrix_r[913*12+:12]), .i_data_2(matrix_i[913*12+:12]), .o_data(c_plus_d[145][3]), .i_clk(i_clk));
Add0000000001  u_0000000397_Add0000000001(.i_data_1(matrix_r[914*12+:12]), .i_data_2(matrix_i[914*12+:12]), .o_data(c_plus_d[146][3]), .i_clk(i_clk));
Add0000000001  u_0000000398_Add0000000001(.i_data_1(matrix_r[915*12+:12]), .i_data_2(matrix_i[915*12+:12]), .o_data(c_plus_d[147][3]), .i_clk(i_clk));
Add0000000001  u_0000000399_Add0000000001(.i_data_1(matrix_r[916*12+:12]), .i_data_2(matrix_i[916*12+:12]), .o_data(c_plus_d[148][3]), .i_clk(i_clk));
Add0000000001  u_000000039A_Add0000000001(.i_data_1(matrix_r[917*12+:12]), .i_data_2(matrix_i[917*12+:12]), .o_data(c_plus_d[149][3]), .i_clk(i_clk));
Add0000000001  u_000000039B_Add0000000001(.i_data_1(matrix_r[918*12+:12]), .i_data_2(matrix_i[918*12+:12]), .o_data(c_plus_d[150][3]), .i_clk(i_clk));
Add0000000001  u_000000039C_Add0000000001(.i_data_1(matrix_r[919*12+:12]), .i_data_2(matrix_i[919*12+:12]), .o_data(c_plus_d[151][3]), .i_clk(i_clk));
Add0000000001  u_000000039D_Add0000000001(.i_data_1(matrix_r[920*12+:12]), .i_data_2(matrix_i[920*12+:12]), .o_data(c_plus_d[152][3]), .i_clk(i_clk));
Add0000000001  u_000000039E_Add0000000001(.i_data_1(matrix_r[921*12+:12]), .i_data_2(matrix_i[921*12+:12]), .o_data(c_plus_d[153][3]), .i_clk(i_clk));
Add0000000001  u_000000039F_Add0000000001(.i_data_1(matrix_r[922*12+:12]), .i_data_2(matrix_i[922*12+:12]), .o_data(c_plus_d[154][3]), .i_clk(i_clk));
Add0000000001  u_00000003A0_Add0000000001(.i_data_1(matrix_r[923*12+:12]), .i_data_2(matrix_i[923*12+:12]), .o_data(c_plus_d[155][3]), .i_clk(i_clk));
Add0000000001  u_00000003A1_Add0000000001(.i_data_1(matrix_r[924*12+:12]), .i_data_2(matrix_i[924*12+:12]), .o_data(c_plus_d[156][3]), .i_clk(i_clk));
Add0000000001  u_00000003A2_Add0000000001(.i_data_1(matrix_r[925*12+:12]), .i_data_2(matrix_i[925*12+:12]), .o_data(c_plus_d[157][3]), .i_clk(i_clk));
Add0000000001  u_00000003A3_Add0000000001(.i_data_1(matrix_r[926*12+:12]), .i_data_2(matrix_i[926*12+:12]), .o_data(c_plus_d[158][3]), .i_clk(i_clk));
Add0000000001  u_00000003A4_Add0000000001(.i_data_1(matrix_r[927*12+:12]), .i_data_2(matrix_i[927*12+:12]), .o_data(c_plus_d[159][3]), .i_clk(i_clk));
Add0000000001  u_00000003A5_Add0000000001(.i_data_1(matrix_r[928*12+:12]), .i_data_2(matrix_i[928*12+:12]), .o_data(c_plus_d[160][3]), .i_clk(i_clk));
Add0000000001  u_00000003A6_Add0000000001(.i_data_1(matrix_r[929*12+:12]), .i_data_2(matrix_i[929*12+:12]), .o_data(c_plus_d[161][3]), .i_clk(i_clk));
Add0000000001  u_00000003A7_Add0000000001(.i_data_1(matrix_r[930*12+:12]), .i_data_2(matrix_i[930*12+:12]), .o_data(c_plus_d[162][3]), .i_clk(i_clk));
Add0000000001  u_00000003A8_Add0000000001(.i_data_1(matrix_r[931*12+:12]), .i_data_2(matrix_i[931*12+:12]), .o_data(c_plus_d[163][3]), .i_clk(i_clk));
Add0000000001  u_00000003A9_Add0000000001(.i_data_1(matrix_r[932*12+:12]), .i_data_2(matrix_i[932*12+:12]), .o_data(c_plus_d[164][3]), .i_clk(i_clk));
Add0000000001  u_00000003AA_Add0000000001(.i_data_1(matrix_r[933*12+:12]), .i_data_2(matrix_i[933*12+:12]), .o_data(c_plus_d[165][3]), .i_clk(i_clk));
Add0000000001  u_00000003AB_Add0000000001(.i_data_1(matrix_r[934*12+:12]), .i_data_2(matrix_i[934*12+:12]), .o_data(c_plus_d[166][3]), .i_clk(i_clk));
Add0000000001  u_00000003AC_Add0000000001(.i_data_1(matrix_r[935*12+:12]), .i_data_2(matrix_i[935*12+:12]), .o_data(c_plus_d[167][3]), .i_clk(i_clk));
Add0000000001  u_00000003AD_Add0000000001(.i_data_1(matrix_r[936*12+:12]), .i_data_2(matrix_i[936*12+:12]), .o_data(c_plus_d[168][3]), .i_clk(i_clk));
Add0000000001  u_00000003AE_Add0000000001(.i_data_1(matrix_r[937*12+:12]), .i_data_2(matrix_i[937*12+:12]), .o_data(c_plus_d[169][3]), .i_clk(i_clk));
Add0000000001  u_00000003AF_Add0000000001(.i_data_1(matrix_r[938*12+:12]), .i_data_2(matrix_i[938*12+:12]), .o_data(c_plus_d[170][3]), .i_clk(i_clk));
Add0000000001  u_00000003B0_Add0000000001(.i_data_1(matrix_r[939*12+:12]), .i_data_2(matrix_i[939*12+:12]), .o_data(c_plus_d[171][3]), .i_clk(i_clk));
Add0000000001  u_00000003B1_Add0000000001(.i_data_1(matrix_r[940*12+:12]), .i_data_2(matrix_i[940*12+:12]), .o_data(c_plus_d[172][3]), .i_clk(i_clk));
Add0000000001  u_00000003B2_Add0000000001(.i_data_1(matrix_r[941*12+:12]), .i_data_2(matrix_i[941*12+:12]), .o_data(c_plus_d[173][3]), .i_clk(i_clk));
Add0000000001  u_00000003B3_Add0000000001(.i_data_1(matrix_r[942*12+:12]), .i_data_2(matrix_i[942*12+:12]), .o_data(c_plus_d[174][3]), .i_clk(i_clk));
Add0000000001  u_00000003B4_Add0000000001(.i_data_1(matrix_r[943*12+:12]), .i_data_2(matrix_i[943*12+:12]), .o_data(c_plus_d[175][3]), .i_clk(i_clk));
Add0000000001  u_00000003B5_Add0000000001(.i_data_1(matrix_r[944*12+:12]), .i_data_2(matrix_i[944*12+:12]), .o_data(c_plus_d[176][3]), .i_clk(i_clk));
Add0000000001  u_00000003B6_Add0000000001(.i_data_1(matrix_r[945*12+:12]), .i_data_2(matrix_i[945*12+:12]), .o_data(c_plus_d[177][3]), .i_clk(i_clk));
Add0000000001  u_00000003B7_Add0000000001(.i_data_1(matrix_r[946*12+:12]), .i_data_2(matrix_i[946*12+:12]), .o_data(c_plus_d[178][3]), .i_clk(i_clk));
Add0000000001  u_00000003B8_Add0000000001(.i_data_1(matrix_r[947*12+:12]), .i_data_2(matrix_i[947*12+:12]), .o_data(c_plus_d[179][3]), .i_clk(i_clk));
Add0000000001  u_00000003B9_Add0000000001(.i_data_1(matrix_r[948*12+:12]), .i_data_2(matrix_i[948*12+:12]), .o_data(c_plus_d[180][3]), .i_clk(i_clk));
Add0000000001  u_00000003BA_Add0000000001(.i_data_1(matrix_r[949*12+:12]), .i_data_2(matrix_i[949*12+:12]), .o_data(c_plus_d[181][3]), .i_clk(i_clk));
Add0000000001  u_00000003BB_Add0000000001(.i_data_1(matrix_r[950*12+:12]), .i_data_2(matrix_i[950*12+:12]), .o_data(c_plus_d[182][3]), .i_clk(i_clk));
Add0000000001  u_00000003BC_Add0000000001(.i_data_1(matrix_r[951*12+:12]), .i_data_2(matrix_i[951*12+:12]), .o_data(c_plus_d[183][3]), .i_clk(i_clk));
Add0000000001  u_00000003BD_Add0000000001(.i_data_1(matrix_r[952*12+:12]), .i_data_2(matrix_i[952*12+:12]), .o_data(c_plus_d[184][3]), .i_clk(i_clk));
Add0000000001  u_00000003BE_Add0000000001(.i_data_1(matrix_r[953*12+:12]), .i_data_2(matrix_i[953*12+:12]), .o_data(c_plus_d[185][3]), .i_clk(i_clk));
Add0000000001  u_00000003BF_Add0000000001(.i_data_1(matrix_r[954*12+:12]), .i_data_2(matrix_i[954*12+:12]), .o_data(c_plus_d[186][3]), .i_clk(i_clk));
Add0000000001  u_00000003C0_Add0000000001(.i_data_1(matrix_r[955*12+:12]), .i_data_2(matrix_i[955*12+:12]), .o_data(c_plus_d[187][3]), .i_clk(i_clk));
Add0000000001  u_00000003C1_Add0000000001(.i_data_1(matrix_r[956*12+:12]), .i_data_2(matrix_i[956*12+:12]), .o_data(c_plus_d[188][3]), .i_clk(i_clk));
Add0000000001  u_00000003C2_Add0000000001(.i_data_1(matrix_r[957*12+:12]), .i_data_2(matrix_i[957*12+:12]), .o_data(c_plus_d[189][3]), .i_clk(i_clk));
Add0000000001  u_00000003C3_Add0000000001(.i_data_1(matrix_r[958*12+:12]), .i_data_2(matrix_i[958*12+:12]), .o_data(c_plus_d[190][3]), .i_clk(i_clk));
Add0000000001  u_00000003C4_Add0000000001(.i_data_1(matrix_r[959*12+:12]), .i_data_2(matrix_i[959*12+:12]), .o_data(c_plus_d[191][3]), .i_clk(i_clk));
Add0000000001  u_00000003C5_Add0000000001(.i_data_1(matrix_r[960*12+:12]), .i_data_2(matrix_i[960*12+:12]), .o_data(c_plus_d[192][3]), .i_clk(i_clk));
Add0000000001  u_00000003C6_Add0000000001(.i_data_1(matrix_r[961*12+:12]), .i_data_2(matrix_i[961*12+:12]), .o_data(c_plus_d[193][3]), .i_clk(i_clk));
Add0000000001  u_00000003C7_Add0000000001(.i_data_1(matrix_r[962*12+:12]), .i_data_2(matrix_i[962*12+:12]), .o_data(c_plus_d[194][3]), .i_clk(i_clk));
Add0000000001  u_00000003C8_Add0000000001(.i_data_1(matrix_r[963*12+:12]), .i_data_2(matrix_i[963*12+:12]), .o_data(c_plus_d[195][3]), .i_clk(i_clk));
Add0000000001  u_00000003C9_Add0000000001(.i_data_1(matrix_r[964*12+:12]), .i_data_2(matrix_i[964*12+:12]), .o_data(c_plus_d[196][3]), .i_clk(i_clk));
Add0000000001  u_00000003CA_Add0000000001(.i_data_1(matrix_r[965*12+:12]), .i_data_2(matrix_i[965*12+:12]), .o_data(c_plus_d[197][3]), .i_clk(i_clk));
Add0000000001  u_00000003CB_Add0000000001(.i_data_1(matrix_r[966*12+:12]), .i_data_2(matrix_i[966*12+:12]), .o_data(c_plus_d[198][3]), .i_clk(i_clk));
Add0000000001  u_00000003CC_Add0000000001(.i_data_1(matrix_r[967*12+:12]), .i_data_2(matrix_i[967*12+:12]), .o_data(c_plus_d[199][3]), .i_clk(i_clk));
Add0000000001  u_00000003CD_Add0000000001(.i_data_1(matrix_r[968*12+:12]), .i_data_2(matrix_i[968*12+:12]), .o_data(c_plus_d[200][3]), .i_clk(i_clk));
Add0000000001  u_00000003CE_Add0000000001(.i_data_1(matrix_r[969*12+:12]), .i_data_2(matrix_i[969*12+:12]), .o_data(c_plus_d[201][3]), .i_clk(i_clk));
Add0000000001  u_00000003CF_Add0000000001(.i_data_1(matrix_r[970*12+:12]), .i_data_2(matrix_i[970*12+:12]), .o_data(c_plus_d[202][3]), .i_clk(i_clk));
Add0000000001  u_00000003D0_Add0000000001(.i_data_1(matrix_r[971*12+:12]), .i_data_2(matrix_i[971*12+:12]), .o_data(c_plus_d[203][3]), .i_clk(i_clk));
Add0000000001  u_00000003D1_Add0000000001(.i_data_1(matrix_r[972*12+:12]), .i_data_2(matrix_i[972*12+:12]), .o_data(c_plus_d[204][3]), .i_clk(i_clk));
Add0000000001  u_00000003D2_Add0000000001(.i_data_1(matrix_r[973*12+:12]), .i_data_2(matrix_i[973*12+:12]), .o_data(c_plus_d[205][3]), .i_clk(i_clk));
Add0000000001  u_00000003D3_Add0000000001(.i_data_1(matrix_r[974*12+:12]), .i_data_2(matrix_i[974*12+:12]), .o_data(c_plus_d[206][3]), .i_clk(i_clk));
Add0000000001  u_00000003D4_Add0000000001(.i_data_1(matrix_r[975*12+:12]), .i_data_2(matrix_i[975*12+:12]), .o_data(c_plus_d[207][3]), .i_clk(i_clk));
Add0000000001  u_00000003D5_Add0000000001(.i_data_1(matrix_r[976*12+:12]), .i_data_2(matrix_i[976*12+:12]), .o_data(c_plus_d[208][3]), .i_clk(i_clk));
Add0000000001  u_00000003D6_Add0000000001(.i_data_1(matrix_r[977*12+:12]), .i_data_2(matrix_i[977*12+:12]), .o_data(c_plus_d[209][3]), .i_clk(i_clk));
Add0000000001  u_00000003D7_Add0000000001(.i_data_1(matrix_r[978*12+:12]), .i_data_2(matrix_i[978*12+:12]), .o_data(c_plus_d[210][3]), .i_clk(i_clk));
Add0000000001  u_00000003D8_Add0000000001(.i_data_1(matrix_r[979*12+:12]), .i_data_2(matrix_i[979*12+:12]), .o_data(c_plus_d[211][3]), .i_clk(i_clk));
Add0000000001  u_00000003D9_Add0000000001(.i_data_1(matrix_r[980*12+:12]), .i_data_2(matrix_i[980*12+:12]), .o_data(c_plus_d[212][3]), .i_clk(i_clk));
Add0000000001  u_00000003DA_Add0000000001(.i_data_1(matrix_r[981*12+:12]), .i_data_2(matrix_i[981*12+:12]), .o_data(c_plus_d[213][3]), .i_clk(i_clk));
Add0000000001  u_00000003DB_Add0000000001(.i_data_1(matrix_r[982*12+:12]), .i_data_2(matrix_i[982*12+:12]), .o_data(c_plus_d[214][3]), .i_clk(i_clk));
Add0000000001  u_00000003DC_Add0000000001(.i_data_1(matrix_r[983*12+:12]), .i_data_2(matrix_i[983*12+:12]), .o_data(c_plus_d[215][3]), .i_clk(i_clk));
Add0000000001  u_00000003DD_Add0000000001(.i_data_1(matrix_r[984*12+:12]), .i_data_2(matrix_i[984*12+:12]), .o_data(c_plus_d[216][3]), .i_clk(i_clk));
Add0000000001  u_00000003DE_Add0000000001(.i_data_1(matrix_r[985*12+:12]), .i_data_2(matrix_i[985*12+:12]), .o_data(c_plus_d[217][3]), .i_clk(i_clk));
Add0000000001  u_00000003DF_Add0000000001(.i_data_1(matrix_r[986*12+:12]), .i_data_2(matrix_i[986*12+:12]), .o_data(c_plus_d[218][3]), .i_clk(i_clk));
Add0000000001  u_00000003E0_Add0000000001(.i_data_1(matrix_r[987*12+:12]), .i_data_2(matrix_i[987*12+:12]), .o_data(c_plus_d[219][3]), .i_clk(i_clk));
Add0000000001  u_00000003E1_Add0000000001(.i_data_1(matrix_r[988*12+:12]), .i_data_2(matrix_i[988*12+:12]), .o_data(c_plus_d[220][3]), .i_clk(i_clk));
Add0000000001  u_00000003E2_Add0000000001(.i_data_1(matrix_r[989*12+:12]), .i_data_2(matrix_i[989*12+:12]), .o_data(c_plus_d[221][3]), .i_clk(i_clk));
Add0000000001  u_00000003E3_Add0000000001(.i_data_1(matrix_r[990*12+:12]), .i_data_2(matrix_i[990*12+:12]), .o_data(c_plus_d[222][3]), .i_clk(i_clk));
Add0000000001  u_00000003E4_Add0000000001(.i_data_1(matrix_r[991*12+:12]), .i_data_2(matrix_i[991*12+:12]), .o_data(c_plus_d[223][3]), .i_clk(i_clk));
Add0000000001  u_00000003E5_Add0000000001(.i_data_1(matrix_r[992*12+:12]), .i_data_2(matrix_i[992*12+:12]), .o_data(c_plus_d[224][3]), .i_clk(i_clk));
Add0000000001  u_00000003E6_Add0000000001(.i_data_1(matrix_r[993*12+:12]), .i_data_2(matrix_i[993*12+:12]), .o_data(c_plus_d[225][3]), .i_clk(i_clk));
Add0000000001  u_00000003E7_Add0000000001(.i_data_1(matrix_r[994*12+:12]), .i_data_2(matrix_i[994*12+:12]), .o_data(c_plus_d[226][3]), .i_clk(i_clk));
Add0000000001  u_00000003E8_Add0000000001(.i_data_1(matrix_r[995*12+:12]), .i_data_2(matrix_i[995*12+:12]), .o_data(c_plus_d[227][3]), .i_clk(i_clk));
Add0000000001  u_00000003E9_Add0000000001(.i_data_1(matrix_r[996*12+:12]), .i_data_2(matrix_i[996*12+:12]), .o_data(c_plus_d[228][3]), .i_clk(i_clk));
Add0000000001  u_00000003EA_Add0000000001(.i_data_1(matrix_r[997*12+:12]), .i_data_2(matrix_i[997*12+:12]), .o_data(c_plus_d[229][3]), .i_clk(i_clk));
Add0000000001  u_00000003EB_Add0000000001(.i_data_1(matrix_r[998*12+:12]), .i_data_2(matrix_i[998*12+:12]), .o_data(c_plus_d[230][3]), .i_clk(i_clk));
Add0000000001  u_00000003EC_Add0000000001(.i_data_1(matrix_r[999*12+:12]), .i_data_2(matrix_i[999*12+:12]), .o_data(c_plus_d[231][3]), .i_clk(i_clk));
Add0000000001  u_00000003ED_Add0000000001(.i_data_1(matrix_r[1000*12+:12]), .i_data_2(matrix_i[1000*12+:12]), .o_data(c_plus_d[232][3]), .i_clk(i_clk));
Add0000000001  u_00000003EE_Add0000000001(.i_data_1(matrix_r[1001*12+:12]), .i_data_2(matrix_i[1001*12+:12]), .o_data(c_plus_d[233][3]), .i_clk(i_clk));
Add0000000001  u_00000003EF_Add0000000001(.i_data_1(matrix_r[1002*12+:12]), .i_data_2(matrix_i[1002*12+:12]), .o_data(c_plus_d[234][3]), .i_clk(i_clk));
Add0000000001  u_00000003F0_Add0000000001(.i_data_1(matrix_r[1003*12+:12]), .i_data_2(matrix_i[1003*12+:12]), .o_data(c_plus_d[235][3]), .i_clk(i_clk));
Add0000000001  u_00000003F1_Add0000000001(.i_data_1(matrix_r[1004*12+:12]), .i_data_2(matrix_i[1004*12+:12]), .o_data(c_plus_d[236][3]), .i_clk(i_clk));
Add0000000001  u_00000003F2_Add0000000001(.i_data_1(matrix_r[1005*12+:12]), .i_data_2(matrix_i[1005*12+:12]), .o_data(c_plus_d[237][3]), .i_clk(i_clk));
Add0000000001  u_00000003F3_Add0000000001(.i_data_1(matrix_r[1006*12+:12]), .i_data_2(matrix_i[1006*12+:12]), .o_data(c_plus_d[238][3]), .i_clk(i_clk));
Add0000000001  u_00000003F4_Add0000000001(.i_data_1(matrix_r[1007*12+:12]), .i_data_2(matrix_i[1007*12+:12]), .o_data(c_plus_d[239][3]), .i_clk(i_clk));
Add0000000001  u_00000003F5_Add0000000001(.i_data_1(matrix_r[1008*12+:12]), .i_data_2(matrix_i[1008*12+:12]), .o_data(c_plus_d[240][3]), .i_clk(i_clk));
Add0000000001  u_00000003F6_Add0000000001(.i_data_1(matrix_r[1009*12+:12]), .i_data_2(matrix_i[1009*12+:12]), .o_data(c_plus_d[241][3]), .i_clk(i_clk));
Add0000000001  u_00000003F7_Add0000000001(.i_data_1(matrix_r[1010*12+:12]), .i_data_2(matrix_i[1010*12+:12]), .o_data(c_plus_d[242][3]), .i_clk(i_clk));
Add0000000001  u_00000003F8_Add0000000001(.i_data_1(matrix_r[1011*12+:12]), .i_data_2(matrix_i[1011*12+:12]), .o_data(c_plus_d[243][3]), .i_clk(i_clk));
Add0000000001  u_00000003F9_Add0000000001(.i_data_1(matrix_r[1012*12+:12]), .i_data_2(matrix_i[1012*12+:12]), .o_data(c_plus_d[244][3]), .i_clk(i_clk));
Add0000000001  u_00000003FA_Add0000000001(.i_data_1(matrix_r[1013*12+:12]), .i_data_2(matrix_i[1013*12+:12]), .o_data(c_plus_d[245][3]), .i_clk(i_clk));
Add0000000001  u_00000003FB_Add0000000001(.i_data_1(matrix_r[1014*12+:12]), .i_data_2(matrix_i[1014*12+:12]), .o_data(c_plus_d[246][3]), .i_clk(i_clk));
Add0000000001  u_00000003FC_Add0000000001(.i_data_1(matrix_r[1015*12+:12]), .i_data_2(matrix_i[1015*12+:12]), .o_data(c_plus_d[247][3]), .i_clk(i_clk));
Add0000000001  u_00000003FD_Add0000000001(.i_data_1(matrix_r[1016*12+:12]), .i_data_2(matrix_i[1016*12+:12]), .o_data(c_plus_d[248][3]), .i_clk(i_clk));
Add0000000001  u_00000003FE_Add0000000001(.i_data_1(matrix_r[1017*12+:12]), .i_data_2(matrix_i[1017*12+:12]), .o_data(c_plus_d[249][3]), .i_clk(i_clk));
Add0000000001  u_00000003FF_Add0000000001(.i_data_1(matrix_r[1018*12+:12]), .i_data_2(matrix_i[1018*12+:12]), .o_data(c_plus_d[250][3]), .i_clk(i_clk));
Add0000000001  u_0000000400_Add0000000001(.i_data_1(matrix_r[1019*12+:12]), .i_data_2(matrix_i[1019*12+:12]), .o_data(c_plus_d[251][3]), .i_clk(i_clk));
Add0000000001  u_0000000401_Add0000000001(.i_data_1(matrix_r[1020*12+:12]), .i_data_2(matrix_i[1020*12+:12]), .o_data(c_plus_d[252][3]), .i_clk(i_clk));
Add0000000001  u_0000000402_Add0000000001(.i_data_1(matrix_r[1021*12+:12]), .i_data_2(matrix_i[1021*12+:12]), .o_data(c_plus_d[253][3]), .i_clk(i_clk));
Add0000000001  u_0000000403_Add0000000001(.i_data_1(matrix_r[1022*12+:12]), .i_data_2(matrix_i[1022*12+:12]), .o_data(c_plus_d[254][3]), .i_clk(i_clk));
Add0000000001  u_0000000404_Add0000000001(.i_data_1(matrix_r[1023*12+:12]), .i_data_2(matrix_i[1023*12+:12]), .o_data(c_plus_d[255][3]), .i_clk(i_clk));
 // L1 Pipeline Registers
 wire [256*4*12-1:0] matrix_r_d, matrix_i_d;
 wire [4*12-1:0] vector_i_d;
Delay0000000005  u_0000000001_Delay0000000005(.i_data(matrix_r), .o_data(matrix_r_d), .i_clk(i_clk));
Delay0000000005  u_0000000002_Delay0000000005(.i_data(matrix_i), .o_data(matrix_i_d), .i_clk(i_clk));
Delay0000000006  u_0000000001_Delay0000000006(.i_data(vector_i), .o_data(vector_i_d), .i_clk(i_clk));
 // Layer 2: Multiply
 wire [12-1:0] A [0:256-1][0:4-1];
 wire [12-1:0] B [0:256-1][0:4-1];
 wire [12-1:0] C [0:256-1][0:4-1];
Mul0000000001  u_0000000001_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[0*12+:12]), .o_data(A[0][0]), .i_clk(i_clk));
Mul0000000001  u_0000000002_Mul0000000001(.i_data_1(c_plus_d[0][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[0][0]), .i_clk(i_clk));
Mul0000000001  u_0000000003_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[0*12+:12]), .o_data(C[0][0]), .i_clk(i_clk));
Mul0000000001  u_0000000004_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[256*12+:12]), .o_data(A[0][1]), .i_clk(i_clk));
Mul0000000001  u_0000000005_Mul0000000001(.i_data_1(c_plus_d[0][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[0][1]), .i_clk(i_clk));
Mul0000000001  u_0000000006_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[256*12+:12]), .o_data(C[0][1]), .i_clk(i_clk));
Mul0000000001  u_0000000007_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[512*12+:12]), .o_data(A[0][2]), .i_clk(i_clk));
Mul0000000001  u_0000000008_Mul0000000001(.i_data_1(c_plus_d[0][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[0][2]), .i_clk(i_clk));
Mul0000000001  u_0000000009_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[512*12+:12]), .o_data(C[0][2]), .i_clk(i_clk));
Mul0000000001  u_000000000A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[768*12+:12]), .o_data(A[0][3]), .i_clk(i_clk));
Mul0000000001  u_000000000B_Mul0000000001(.i_data_1(c_plus_d[0][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[0][3]), .i_clk(i_clk));
Mul0000000001  u_000000000C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[768*12+:12]), .o_data(C[0][3]), .i_clk(i_clk));
Mul0000000001  u_000000000D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[1*12+:12]), .o_data(A[1][0]), .i_clk(i_clk));
Mul0000000001  u_000000000E_Mul0000000001(.i_data_1(c_plus_d[1][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[1][0]), .i_clk(i_clk));
Mul0000000001  u_000000000F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[1*12+:12]), .o_data(C[1][0]), .i_clk(i_clk));
Mul0000000001  u_0000000010_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[257*12+:12]), .o_data(A[1][1]), .i_clk(i_clk));
Mul0000000001  u_0000000011_Mul0000000001(.i_data_1(c_plus_d[1][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[1][1]), .i_clk(i_clk));
Mul0000000001  u_0000000012_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[257*12+:12]), .o_data(C[1][1]), .i_clk(i_clk));
Mul0000000001  u_0000000013_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[513*12+:12]), .o_data(A[1][2]), .i_clk(i_clk));
Mul0000000001  u_0000000014_Mul0000000001(.i_data_1(c_plus_d[1][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[1][2]), .i_clk(i_clk));
Mul0000000001  u_0000000015_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[513*12+:12]), .o_data(C[1][2]), .i_clk(i_clk));
Mul0000000001  u_0000000016_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[769*12+:12]), .o_data(A[1][3]), .i_clk(i_clk));
Mul0000000001  u_0000000017_Mul0000000001(.i_data_1(c_plus_d[1][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[1][3]), .i_clk(i_clk));
Mul0000000001  u_0000000018_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[769*12+:12]), .o_data(C[1][3]), .i_clk(i_clk));
Mul0000000001  u_0000000019_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[2*12+:12]), .o_data(A[2][0]), .i_clk(i_clk));
Mul0000000001  u_000000001A_Mul0000000001(.i_data_1(c_plus_d[2][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[2][0]), .i_clk(i_clk));
Mul0000000001  u_000000001B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[2*12+:12]), .o_data(C[2][0]), .i_clk(i_clk));
Mul0000000001  u_000000001C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[258*12+:12]), .o_data(A[2][1]), .i_clk(i_clk));
Mul0000000001  u_000000001D_Mul0000000001(.i_data_1(c_plus_d[2][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[2][1]), .i_clk(i_clk));
Mul0000000001  u_000000001E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[258*12+:12]), .o_data(C[2][1]), .i_clk(i_clk));
Mul0000000001  u_000000001F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[514*12+:12]), .o_data(A[2][2]), .i_clk(i_clk));
Mul0000000001  u_0000000020_Mul0000000001(.i_data_1(c_plus_d[2][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[2][2]), .i_clk(i_clk));
Mul0000000001  u_0000000021_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[514*12+:12]), .o_data(C[2][2]), .i_clk(i_clk));
Mul0000000001  u_0000000022_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[770*12+:12]), .o_data(A[2][3]), .i_clk(i_clk));
Mul0000000001  u_0000000023_Mul0000000001(.i_data_1(c_plus_d[2][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[2][3]), .i_clk(i_clk));
Mul0000000001  u_0000000024_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[770*12+:12]), .o_data(C[2][3]), .i_clk(i_clk));
Mul0000000001  u_0000000025_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[3*12+:12]), .o_data(A[3][0]), .i_clk(i_clk));
Mul0000000001  u_0000000026_Mul0000000001(.i_data_1(c_plus_d[3][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[3][0]), .i_clk(i_clk));
Mul0000000001  u_0000000027_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[3*12+:12]), .o_data(C[3][0]), .i_clk(i_clk));
Mul0000000001  u_0000000028_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[259*12+:12]), .o_data(A[3][1]), .i_clk(i_clk));
Mul0000000001  u_0000000029_Mul0000000001(.i_data_1(c_plus_d[3][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[3][1]), .i_clk(i_clk));
Mul0000000001  u_000000002A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[259*12+:12]), .o_data(C[3][1]), .i_clk(i_clk));
Mul0000000001  u_000000002B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[515*12+:12]), .o_data(A[3][2]), .i_clk(i_clk));
Mul0000000001  u_000000002C_Mul0000000001(.i_data_1(c_plus_d[3][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[3][2]), .i_clk(i_clk));
Mul0000000001  u_000000002D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[515*12+:12]), .o_data(C[3][2]), .i_clk(i_clk));
Mul0000000001  u_000000002E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[771*12+:12]), .o_data(A[3][3]), .i_clk(i_clk));
Mul0000000001  u_000000002F_Mul0000000001(.i_data_1(c_plus_d[3][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[3][3]), .i_clk(i_clk));
Mul0000000001  u_0000000030_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[771*12+:12]), .o_data(C[3][3]), .i_clk(i_clk));
Mul0000000001  u_0000000031_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[4*12+:12]), .o_data(A[4][0]), .i_clk(i_clk));
Mul0000000001  u_0000000032_Mul0000000001(.i_data_1(c_plus_d[4][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[4][0]), .i_clk(i_clk));
Mul0000000001  u_0000000033_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[4*12+:12]), .o_data(C[4][0]), .i_clk(i_clk));
Mul0000000001  u_0000000034_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[260*12+:12]), .o_data(A[4][1]), .i_clk(i_clk));
Mul0000000001  u_0000000035_Mul0000000001(.i_data_1(c_plus_d[4][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[4][1]), .i_clk(i_clk));
Mul0000000001  u_0000000036_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[260*12+:12]), .o_data(C[4][1]), .i_clk(i_clk));
Mul0000000001  u_0000000037_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[516*12+:12]), .o_data(A[4][2]), .i_clk(i_clk));
Mul0000000001  u_0000000038_Mul0000000001(.i_data_1(c_plus_d[4][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[4][2]), .i_clk(i_clk));
Mul0000000001  u_0000000039_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[516*12+:12]), .o_data(C[4][2]), .i_clk(i_clk));
Mul0000000001  u_000000003A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[772*12+:12]), .o_data(A[4][3]), .i_clk(i_clk));
Mul0000000001  u_000000003B_Mul0000000001(.i_data_1(c_plus_d[4][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[4][3]), .i_clk(i_clk));
Mul0000000001  u_000000003C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[772*12+:12]), .o_data(C[4][3]), .i_clk(i_clk));
Mul0000000001  u_000000003D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[5*12+:12]), .o_data(A[5][0]), .i_clk(i_clk));
Mul0000000001  u_000000003E_Mul0000000001(.i_data_1(c_plus_d[5][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[5][0]), .i_clk(i_clk));
Mul0000000001  u_000000003F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[5*12+:12]), .o_data(C[5][0]), .i_clk(i_clk));
Mul0000000001  u_0000000040_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[261*12+:12]), .o_data(A[5][1]), .i_clk(i_clk));
Mul0000000001  u_0000000041_Mul0000000001(.i_data_1(c_plus_d[5][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[5][1]), .i_clk(i_clk));
Mul0000000001  u_0000000042_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[261*12+:12]), .o_data(C[5][1]), .i_clk(i_clk));
Mul0000000001  u_0000000043_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[517*12+:12]), .o_data(A[5][2]), .i_clk(i_clk));
Mul0000000001  u_0000000044_Mul0000000001(.i_data_1(c_plus_d[5][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[5][2]), .i_clk(i_clk));
Mul0000000001  u_0000000045_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[517*12+:12]), .o_data(C[5][2]), .i_clk(i_clk));
Mul0000000001  u_0000000046_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[773*12+:12]), .o_data(A[5][3]), .i_clk(i_clk));
Mul0000000001  u_0000000047_Mul0000000001(.i_data_1(c_plus_d[5][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[5][3]), .i_clk(i_clk));
Mul0000000001  u_0000000048_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[773*12+:12]), .o_data(C[5][3]), .i_clk(i_clk));
Mul0000000001  u_0000000049_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[6*12+:12]), .o_data(A[6][0]), .i_clk(i_clk));
Mul0000000001  u_000000004A_Mul0000000001(.i_data_1(c_plus_d[6][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[6][0]), .i_clk(i_clk));
Mul0000000001  u_000000004B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[6*12+:12]), .o_data(C[6][0]), .i_clk(i_clk));
Mul0000000001  u_000000004C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[262*12+:12]), .o_data(A[6][1]), .i_clk(i_clk));
Mul0000000001  u_000000004D_Mul0000000001(.i_data_1(c_plus_d[6][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[6][1]), .i_clk(i_clk));
Mul0000000001  u_000000004E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[262*12+:12]), .o_data(C[6][1]), .i_clk(i_clk));
Mul0000000001  u_000000004F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[518*12+:12]), .o_data(A[6][2]), .i_clk(i_clk));
Mul0000000001  u_0000000050_Mul0000000001(.i_data_1(c_plus_d[6][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[6][2]), .i_clk(i_clk));
Mul0000000001  u_0000000051_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[518*12+:12]), .o_data(C[6][2]), .i_clk(i_clk));
Mul0000000001  u_0000000052_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[774*12+:12]), .o_data(A[6][3]), .i_clk(i_clk));
Mul0000000001  u_0000000053_Mul0000000001(.i_data_1(c_plus_d[6][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[6][3]), .i_clk(i_clk));
Mul0000000001  u_0000000054_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[774*12+:12]), .o_data(C[6][3]), .i_clk(i_clk));
Mul0000000001  u_0000000055_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[7*12+:12]), .o_data(A[7][0]), .i_clk(i_clk));
Mul0000000001  u_0000000056_Mul0000000001(.i_data_1(c_plus_d[7][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[7][0]), .i_clk(i_clk));
Mul0000000001  u_0000000057_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[7*12+:12]), .o_data(C[7][0]), .i_clk(i_clk));
Mul0000000001  u_0000000058_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[263*12+:12]), .o_data(A[7][1]), .i_clk(i_clk));
Mul0000000001  u_0000000059_Mul0000000001(.i_data_1(c_plus_d[7][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[7][1]), .i_clk(i_clk));
Mul0000000001  u_000000005A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[263*12+:12]), .o_data(C[7][1]), .i_clk(i_clk));
Mul0000000001  u_000000005B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[519*12+:12]), .o_data(A[7][2]), .i_clk(i_clk));
Mul0000000001  u_000000005C_Mul0000000001(.i_data_1(c_plus_d[7][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[7][2]), .i_clk(i_clk));
Mul0000000001  u_000000005D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[519*12+:12]), .o_data(C[7][2]), .i_clk(i_clk));
Mul0000000001  u_000000005E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[775*12+:12]), .o_data(A[7][3]), .i_clk(i_clk));
Mul0000000001  u_000000005F_Mul0000000001(.i_data_1(c_plus_d[7][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[7][3]), .i_clk(i_clk));
Mul0000000001  u_0000000060_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[775*12+:12]), .o_data(C[7][3]), .i_clk(i_clk));
Mul0000000001  u_0000000061_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[8*12+:12]), .o_data(A[8][0]), .i_clk(i_clk));
Mul0000000001  u_0000000062_Mul0000000001(.i_data_1(c_plus_d[8][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[8][0]), .i_clk(i_clk));
Mul0000000001  u_0000000063_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[8*12+:12]), .o_data(C[8][0]), .i_clk(i_clk));
Mul0000000001  u_0000000064_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[264*12+:12]), .o_data(A[8][1]), .i_clk(i_clk));
Mul0000000001  u_0000000065_Mul0000000001(.i_data_1(c_plus_d[8][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[8][1]), .i_clk(i_clk));
Mul0000000001  u_0000000066_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[264*12+:12]), .o_data(C[8][1]), .i_clk(i_clk));
Mul0000000001  u_0000000067_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[520*12+:12]), .o_data(A[8][2]), .i_clk(i_clk));
Mul0000000001  u_0000000068_Mul0000000001(.i_data_1(c_plus_d[8][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[8][2]), .i_clk(i_clk));
Mul0000000001  u_0000000069_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[520*12+:12]), .o_data(C[8][2]), .i_clk(i_clk));
Mul0000000001  u_000000006A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[776*12+:12]), .o_data(A[8][3]), .i_clk(i_clk));
Mul0000000001  u_000000006B_Mul0000000001(.i_data_1(c_plus_d[8][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[8][3]), .i_clk(i_clk));
Mul0000000001  u_000000006C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[776*12+:12]), .o_data(C[8][3]), .i_clk(i_clk));
Mul0000000001  u_000000006D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[9*12+:12]), .o_data(A[9][0]), .i_clk(i_clk));
Mul0000000001  u_000000006E_Mul0000000001(.i_data_1(c_plus_d[9][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[9][0]), .i_clk(i_clk));
Mul0000000001  u_000000006F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[9*12+:12]), .o_data(C[9][0]), .i_clk(i_clk));
Mul0000000001  u_0000000070_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[265*12+:12]), .o_data(A[9][1]), .i_clk(i_clk));
Mul0000000001  u_0000000071_Mul0000000001(.i_data_1(c_plus_d[9][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[9][1]), .i_clk(i_clk));
Mul0000000001  u_0000000072_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[265*12+:12]), .o_data(C[9][1]), .i_clk(i_clk));
Mul0000000001  u_0000000073_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[521*12+:12]), .o_data(A[9][2]), .i_clk(i_clk));
Mul0000000001  u_0000000074_Mul0000000001(.i_data_1(c_plus_d[9][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[9][2]), .i_clk(i_clk));
Mul0000000001  u_0000000075_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[521*12+:12]), .o_data(C[9][2]), .i_clk(i_clk));
Mul0000000001  u_0000000076_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[777*12+:12]), .o_data(A[9][3]), .i_clk(i_clk));
Mul0000000001  u_0000000077_Mul0000000001(.i_data_1(c_plus_d[9][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[9][3]), .i_clk(i_clk));
Mul0000000001  u_0000000078_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[777*12+:12]), .o_data(C[9][3]), .i_clk(i_clk));
Mul0000000001  u_0000000079_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[10*12+:12]), .o_data(A[10][0]), .i_clk(i_clk));
Mul0000000001  u_000000007A_Mul0000000001(.i_data_1(c_plus_d[10][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[10][0]), .i_clk(i_clk));
Mul0000000001  u_000000007B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[10*12+:12]), .o_data(C[10][0]), .i_clk(i_clk));
Mul0000000001  u_000000007C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[266*12+:12]), .o_data(A[10][1]), .i_clk(i_clk));
Mul0000000001  u_000000007D_Mul0000000001(.i_data_1(c_plus_d[10][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[10][1]), .i_clk(i_clk));
Mul0000000001  u_000000007E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[266*12+:12]), .o_data(C[10][1]), .i_clk(i_clk));
Mul0000000001  u_000000007F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[522*12+:12]), .o_data(A[10][2]), .i_clk(i_clk));
Mul0000000001  u_0000000080_Mul0000000001(.i_data_1(c_plus_d[10][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[10][2]), .i_clk(i_clk));
Mul0000000001  u_0000000081_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[522*12+:12]), .o_data(C[10][2]), .i_clk(i_clk));
Mul0000000001  u_0000000082_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[778*12+:12]), .o_data(A[10][3]), .i_clk(i_clk));
Mul0000000001  u_0000000083_Mul0000000001(.i_data_1(c_plus_d[10][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[10][3]), .i_clk(i_clk));
Mul0000000001  u_0000000084_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[778*12+:12]), .o_data(C[10][3]), .i_clk(i_clk));
Mul0000000001  u_0000000085_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[11*12+:12]), .o_data(A[11][0]), .i_clk(i_clk));
Mul0000000001  u_0000000086_Mul0000000001(.i_data_1(c_plus_d[11][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[11][0]), .i_clk(i_clk));
Mul0000000001  u_0000000087_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[11*12+:12]), .o_data(C[11][0]), .i_clk(i_clk));
Mul0000000001  u_0000000088_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[267*12+:12]), .o_data(A[11][1]), .i_clk(i_clk));
Mul0000000001  u_0000000089_Mul0000000001(.i_data_1(c_plus_d[11][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[11][1]), .i_clk(i_clk));
Mul0000000001  u_000000008A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[267*12+:12]), .o_data(C[11][1]), .i_clk(i_clk));
Mul0000000001  u_000000008B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[523*12+:12]), .o_data(A[11][2]), .i_clk(i_clk));
Mul0000000001  u_000000008C_Mul0000000001(.i_data_1(c_plus_d[11][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[11][2]), .i_clk(i_clk));
Mul0000000001  u_000000008D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[523*12+:12]), .o_data(C[11][2]), .i_clk(i_clk));
Mul0000000001  u_000000008E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[779*12+:12]), .o_data(A[11][3]), .i_clk(i_clk));
Mul0000000001  u_000000008F_Mul0000000001(.i_data_1(c_plus_d[11][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[11][3]), .i_clk(i_clk));
Mul0000000001  u_0000000090_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[779*12+:12]), .o_data(C[11][3]), .i_clk(i_clk));
Mul0000000001  u_0000000091_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[12*12+:12]), .o_data(A[12][0]), .i_clk(i_clk));
Mul0000000001  u_0000000092_Mul0000000001(.i_data_1(c_plus_d[12][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[12][0]), .i_clk(i_clk));
Mul0000000001  u_0000000093_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[12*12+:12]), .o_data(C[12][0]), .i_clk(i_clk));
Mul0000000001  u_0000000094_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[268*12+:12]), .o_data(A[12][1]), .i_clk(i_clk));
Mul0000000001  u_0000000095_Mul0000000001(.i_data_1(c_plus_d[12][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[12][1]), .i_clk(i_clk));
Mul0000000001  u_0000000096_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[268*12+:12]), .o_data(C[12][1]), .i_clk(i_clk));
Mul0000000001  u_0000000097_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[524*12+:12]), .o_data(A[12][2]), .i_clk(i_clk));
Mul0000000001  u_0000000098_Mul0000000001(.i_data_1(c_plus_d[12][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[12][2]), .i_clk(i_clk));
Mul0000000001  u_0000000099_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[524*12+:12]), .o_data(C[12][2]), .i_clk(i_clk));
Mul0000000001  u_000000009A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[780*12+:12]), .o_data(A[12][3]), .i_clk(i_clk));
Mul0000000001  u_000000009B_Mul0000000001(.i_data_1(c_plus_d[12][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[12][3]), .i_clk(i_clk));
Mul0000000001  u_000000009C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[780*12+:12]), .o_data(C[12][3]), .i_clk(i_clk));
Mul0000000001  u_000000009D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[13*12+:12]), .o_data(A[13][0]), .i_clk(i_clk));
Mul0000000001  u_000000009E_Mul0000000001(.i_data_1(c_plus_d[13][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[13][0]), .i_clk(i_clk));
Mul0000000001  u_000000009F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[13*12+:12]), .o_data(C[13][0]), .i_clk(i_clk));
Mul0000000001  u_00000000A0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[269*12+:12]), .o_data(A[13][1]), .i_clk(i_clk));
Mul0000000001  u_00000000A1_Mul0000000001(.i_data_1(c_plus_d[13][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[13][1]), .i_clk(i_clk));
Mul0000000001  u_00000000A2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[269*12+:12]), .o_data(C[13][1]), .i_clk(i_clk));
Mul0000000001  u_00000000A3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[525*12+:12]), .o_data(A[13][2]), .i_clk(i_clk));
Mul0000000001  u_00000000A4_Mul0000000001(.i_data_1(c_plus_d[13][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[13][2]), .i_clk(i_clk));
Mul0000000001  u_00000000A5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[525*12+:12]), .o_data(C[13][2]), .i_clk(i_clk));
Mul0000000001  u_00000000A6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[781*12+:12]), .o_data(A[13][3]), .i_clk(i_clk));
Mul0000000001  u_00000000A7_Mul0000000001(.i_data_1(c_plus_d[13][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[13][3]), .i_clk(i_clk));
Mul0000000001  u_00000000A8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[781*12+:12]), .o_data(C[13][3]), .i_clk(i_clk));
Mul0000000001  u_00000000A9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[14*12+:12]), .o_data(A[14][0]), .i_clk(i_clk));
Mul0000000001  u_00000000AA_Mul0000000001(.i_data_1(c_plus_d[14][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[14][0]), .i_clk(i_clk));
Mul0000000001  u_00000000AB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[14*12+:12]), .o_data(C[14][0]), .i_clk(i_clk));
Mul0000000001  u_00000000AC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[270*12+:12]), .o_data(A[14][1]), .i_clk(i_clk));
Mul0000000001  u_00000000AD_Mul0000000001(.i_data_1(c_plus_d[14][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[14][1]), .i_clk(i_clk));
Mul0000000001  u_00000000AE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[270*12+:12]), .o_data(C[14][1]), .i_clk(i_clk));
Mul0000000001  u_00000000AF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[526*12+:12]), .o_data(A[14][2]), .i_clk(i_clk));
Mul0000000001  u_00000000B0_Mul0000000001(.i_data_1(c_plus_d[14][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[14][2]), .i_clk(i_clk));
Mul0000000001  u_00000000B1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[526*12+:12]), .o_data(C[14][2]), .i_clk(i_clk));
Mul0000000001  u_00000000B2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[782*12+:12]), .o_data(A[14][3]), .i_clk(i_clk));
Mul0000000001  u_00000000B3_Mul0000000001(.i_data_1(c_plus_d[14][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[14][3]), .i_clk(i_clk));
Mul0000000001  u_00000000B4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[782*12+:12]), .o_data(C[14][3]), .i_clk(i_clk));
Mul0000000001  u_00000000B5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[15*12+:12]), .o_data(A[15][0]), .i_clk(i_clk));
Mul0000000001  u_00000000B6_Mul0000000001(.i_data_1(c_plus_d[15][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[15][0]), .i_clk(i_clk));
Mul0000000001  u_00000000B7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[15*12+:12]), .o_data(C[15][0]), .i_clk(i_clk));
Mul0000000001  u_00000000B8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[271*12+:12]), .o_data(A[15][1]), .i_clk(i_clk));
Mul0000000001  u_00000000B9_Mul0000000001(.i_data_1(c_plus_d[15][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[15][1]), .i_clk(i_clk));
Mul0000000001  u_00000000BA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[271*12+:12]), .o_data(C[15][1]), .i_clk(i_clk));
Mul0000000001  u_00000000BB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[527*12+:12]), .o_data(A[15][2]), .i_clk(i_clk));
Mul0000000001  u_00000000BC_Mul0000000001(.i_data_1(c_plus_d[15][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[15][2]), .i_clk(i_clk));
Mul0000000001  u_00000000BD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[527*12+:12]), .o_data(C[15][2]), .i_clk(i_clk));
Mul0000000001  u_00000000BE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[783*12+:12]), .o_data(A[15][3]), .i_clk(i_clk));
Mul0000000001  u_00000000BF_Mul0000000001(.i_data_1(c_plus_d[15][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[15][3]), .i_clk(i_clk));
Mul0000000001  u_00000000C0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[783*12+:12]), .o_data(C[15][3]), .i_clk(i_clk));
Mul0000000001  u_00000000C1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[16*12+:12]), .o_data(A[16][0]), .i_clk(i_clk));
Mul0000000001  u_00000000C2_Mul0000000001(.i_data_1(c_plus_d[16][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[16][0]), .i_clk(i_clk));
Mul0000000001  u_00000000C3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[16*12+:12]), .o_data(C[16][0]), .i_clk(i_clk));
Mul0000000001  u_00000000C4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[272*12+:12]), .o_data(A[16][1]), .i_clk(i_clk));
Mul0000000001  u_00000000C5_Mul0000000001(.i_data_1(c_plus_d[16][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[16][1]), .i_clk(i_clk));
Mul0000000001  u_00000000C6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[272*12+:12]), .o_data(C[16][1]), .i_clk(i_clk));
Mul0000000001  u_00000000C7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[528*12+:12]), .o_data(A[16][2]), .i_clk(i_clk));
Mul0000000001  u_00000000C8_Mul0000000001(.i_data_1(c_plus_d[16][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[16][2]), .i_clk(i_clk));
Mul0000000001  u_00000000C9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[528*12+:12]), .o_data(C[16][2]), .i_clk(i_clk));
Mul0000000001  u_00000000CA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[784*12+:12]), .o_data(A[16][3]), .i_clk(i_clk));
Mul0000000001  u_00000000CB_Mul0000000001(.i_data_1(c_plus_d[16][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[16][3]), .i_clk(i_clk));
Mul0000000001  u_00000000CC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[784*12+:12]), .o_data(C[16][3]), .i_clk(i_clk));
Mul0000000001  u_00000000CD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[17*12+:12]), .o_data(A[17][0]), .i_clk(i_clk));
Mul0000000001  u_00000000CE_Mul0000000001(.i_data_1(c_plus_d[17][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[17][0]), .i_clk(i_clk));
Mul0000000001  u_00000000CF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[17*12+:12]), .o_data(C[17][0]), .i_clk(i_clk));
Mul0000000001  u_00000000D0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[273*12+:12]), .o_data(A[17][1]), .i_clk(i_clk));
Mul0000000001  u_00000000D1_Mul0000000001(.i_data_1(c_plus_d[17][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[17][1]), .i_clk(i_clk));
Mul0000000001  u_00000000D2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[273*12+:12]), .o_data(C[17][1]), .i_clk(i_clk));
Mul0000000001  u_00000000D3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[529*12+:12]), .o_data(A[17][2]), .i_clk(i_clk));
Mul0000000001  u_00000000D4_Mul0000000001(.i_data_1(c_plus_d[17][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[17][2]), .i_clk(i_clk));
Mul0000000001  u_00000000D5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[529*12+:12]), .o_data(C[17][2]), .i_clk(i_clk));
Mul0000000001  u_00000000D6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[785*12+:12]), .o_data(A[17][3]), .i_clk(i_clk));
Mul0000000001  u_00000000D7_Mul0000000001(.i_data_1(c_plus_d[17][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[17][3]), .i_clk(i_clk));
Mul0000000001  u_00000000D8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[785*12+:12]), .o_data(C[17][3]), .i_clk(i_clk));
Mul0000000001  u_00000000D9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[18*12+:12]), .o_data(A[18][0]), .i_clk(i_clk));
Mul0000000001  u_00000000DA_Mul0000000001(.i_data_1(c_plus_d[18][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[18][0]), .i_clk(i_clk));
Mul0000000001  u_00000000DB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[18*12+:12]), .o_data(C[18][0]), .i_clk(i_clk));
Mul0000000001  u_00000000DC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[274*12+:12]), .o_data(A[18][1]), .i_clk(i_clk));
Mul0000000001  u_00000000DD_Mul0000000001(.i_data_1(c_plus_d[18][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[18][1]), .i_clk(i_clk));
Mul0000000001  u_00000000DE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[274*12+:12]), .o_data(C[18][1]), .i_clk(i_clk));
Mul0000000001  u_00000000DF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[530*12+:12]), .o_data(A[18][2]), .i_clk(i_clk));
Mul0000000001  u_00000000E0_Mul0000000001(.i_data_1(c_plus_d[18][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[18][2]), .i_clk(i_clk));
Mul0000000001  u_00000000E1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[530*12+:12]), .o_data(C[18][2]), .i_clk(i_clk));
Mul0000000001  u_00000000E2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[786*12+:12]), .o_data(A[18][3]), .i_clk(i_clk));
Mul0000000001  u_00000000E3_Mul0000000001(.i_data_1(c_plus_d[18][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[18][3]), .i_clk(i_clk));
Mul0000000001  u_00000000E4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[786*12+:12]), .o_data(C[18][3]), .i_clk(i_clk));
Mul0000000001  u_00000000E5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[19*12+:12]), .o_data(A[19][0]), .i_clk(i_clk));
Mul0000000001  u_00000000E6_Mul0000000001(.i_data_1(c_plus_d[19][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[19][0]), .i_clk(i_clk));
Mul0000000001  u_00000000E7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[19*12+:12]), .o_data(C[19][0]), .i_clk(i_clk));
Mul0000000001  u_00000000E8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[275*12+:12]), .o_data(A[19][1]), .i_clk(i_clk));
Mul0000000001  u_00000000E9_Mul0000000001(.i_data_1(c_plus_d[19][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[19][1]), .i_clk(i_clk));
Mul0000000001  u_00000000EA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[275*12+:12]), .o_data(C[19][1]), .i_clk(i_clk));
Mul0000000001  u_00000000EB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[531*12+:12]), .o_data(A[19][2]), .i_clk(i_clk));
Mul0000000001  u_00000000EC_Mul0000000001(.i_data_1(c_plus_d[19][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[19][2]), .i_clk(i_clk));
Mul0000000001  u_00000000ED_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[531*12+:12]), .o_data(C[19][2]), .i_clk(i_clk));
Mul0000000001  u_00000000EE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[787*12+:12]), .o_data(A[19][3]), .i_clk(i_clk));
Mul0000000001  u_00000000EF_Mul0000000001(.i_data_1(c_plus_d[19][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[19][3]), .i_clk(i_clk));
Mul0000000001  u_00000000F0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[787*12+:12]), .o_data(C[19][3]), .i_clk(i_clk));
Mul0000000001  u_00000000F1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[20*12+:12]), .o_data(A[20][0]), .i_clk(i_clk));
Mul0000000001  u_00000000F2_Mul0000000001(.i_data_1(c_plus_d[20][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[20][0]), .i_clk(i_clk));
Mul0000000001  u_00000000F3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[20*12+:12]), .o_data(C[20][0]), .i_clk(i_clk));
Mul0000000001  u_00000000F4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[276*12+:12]), .o_data(A[20][1]), .i_clk(i_clk));
Mul0000000001  u_00000000F5_Mul0000000001(.i_data_1(c_plus_d[20][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[20][1]), .i_clk(i_clk));
Mul0000000001  u_00000000F6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[276*12+:12]), .o_data(C[20][1]), .i_clk(i_clk));
Mul0000000001  u_00000000F7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[532*12+:12]), .o_data(A[20][2]), .i_clk(i_clk));
Mul0000000001  u_00000000F8_Mul0000000001(.i_data_1(c_plus_d[20][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[20][2]), .i_clk(i_clk));
Mul0000000001  u_00000000F9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[532*12+:12]), .o_data(C[20][2]), .i_clk(i_clk));
Mul0000000001  u_00000000FA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[788*12+:12]), .o_data(A[20][3]), .i_clk(i_clk));
Mul0000000001  u_00000000FB_Mul0000000001(.i_data_1(c_plus_d[20][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[20][3]), .i_clk(i_clk));
Mul0000000001  u_00000000FC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[788*12+:12]), .o_data(C[20][3]), .i_clk(i_clk));
Mul0000000001  u_00000000FD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[21*12+:12]), .o_data(A[21][0]), .i_clk(i_clk));
Mul0000000001  u_00000000FE_Mul0000000001(.i_data_1(c_plus_d[21][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[21][0]), .i_clk(i_clk));
Mul0000000001  u_00000000FF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[21*12+:12]), .o_data(C[21][0]), .i_clk(i_clk));
Mul0000000001  u_0000000100_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[277*12+:12]), .o_data(A[21][1]), .i_clk(i_clk));
Mul0000000001  u_0000000101_Mul0000000001(.i_data_1(c_plus_d[21][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[21][1]), .i_clk(i_clk));
Mul0000000001  u_0000000102_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[277*12+:12]), .o_data(C[21][1]), .i_clk(i_clk));
Mul0000000001  u_0000000103_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[533*12+:12]), .o_data(A[21][2]), .i_clk(i_clk));
Mul0000000001  u_0000000104_Mul0000000001(.i_data_1(c_plus_d[21][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[21][2]), .i_clk(i_clk));
Mul0000000001  u_0000000105_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[533*12+:12]), .o_data(C[21][2]), .i_clk(i_clk));
Mul0000000001  u_0000000106_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[789*12+:12]), .o_data(A[21][3]), .i_clk(i_clk));
Mul0000000001  u_0000000107_Mul0000000001(.i_data_1(c_plus_d[21][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[21][3]), .i_clk(i_clk));
Mul0000000001  u_0000000108_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[789*12+:12]), .o_data(C[21][3]), .i_clk(i_clk));
Mul0000000001  u_0000000109_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[22*12+:12]), .o_data(A[22][0]), .i_clk(i_clk));
Mul0000000001  u_000000010A_Mul0000000001(.i_data_1(c_plus_d[22][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[22][0]), .i_clk(i_clk));
Mul0000000001  u_000000010B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[22*12+:12]), .o_data(C[22][0]), .i_clk(i_clk));
Mul0000000001  u_000000010C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[278*12+:12]), .o_data(A[22][1]), .i_clk(i_clk));
Mul0000000001  u_000000010D_Mul0000000001(.i_data_1(c_plus_d[22][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[22][1]), .i_clk(i_clk));
Mul0000000001  u_000000010E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[278*12+:12]), .o_data(C[22][1]), .i_clk(i_clk));
Mul0000000001  u_000000010F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[534*12+:12]), .o_data(A[22][2]), .i_clk(i_clk));
Mul0000000001  u_0000000110_Mul0000000001(.i_data_1(c_plus_d[22][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[22][2]), .i_clk(i_clk));
Mul0000000001  u_0000000111_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[534*12+:12]), .o_data(C[22][2]), .i_clk(i_clk));
Mul0000000001  u_0000000112_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[790*12+:12]), .o_data(A[22][3]), .i_clk(i_clk));
Mul0000000001  u_0000000113_Mul0000000001(.i_data_1(c_plus_d[22][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[22][3]), .i_clk(i_clk));
Mul0000000001  u_0000000114_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[790*12+:12]), .o_data(C[22][3]), .i_clk(i_clk));
Mul0000000001  u_0000000115_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[23*12+:12]), .o_data(A[23][0]), .i_clk(i_clk));
Mul0000000001  u_0000000116_Mul0000000001(.i_data_1(c_plus_d[23][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[23][0]), .i_clk(i_clk));
Mul0000000001  u_0000000117_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[23*12+:12]), .o_data(C[23][0]), .i_clk(i_clk));
Mul0000000001  u_0000000118_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[279*12+:12]), .o_data(A[23][1]), .i_clk(i_clk));
Mul0000000001  u_0000000119_Mul0000000001(.i_data_1(c_plus_d[23][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[23][1]), .i_clk(i_clk));
Mul0000000001  u_000000011A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[279*12+:12]), .o_data(C[23][1]), .i_clk(i_clk));
Mul0000000001  u_000000011B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[535*12+:12]), .o_data(A[23][2]), .i_clk(i_clk));
Mul0000000001  u_000000011C_Mul0000000001(.i_data_1(c_plus_d[23][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[23][2]), .i_clk(i_clk));
Mul0000000001  u_000000011D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[535*12+:12]), .o_data(C[23][2]), .i_clk(i_clk));
Mul0000000001  u_000000011E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[791*12+:12]), .o_data(A[23][3]), .i_clk(i_clk));
Mul0000000001  u_000000011F_Mul0000000001(.i_data_1(c_plus_d[23][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[23][3]), .i_clk(i_clk));
Mul0000000001  u_0000000120_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[791*12+:12]), .o_data(C[23][3]), .i_clk(i_clk));
Mul0000000001  u_0000000121_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[24*12+:12]), .o_data(A[24][0]), .i_clk(i_clk));
Mul0000000001  u_0000000122_Mul0000000001(.i_data_1(c_plus_d[24][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[24][0]), .i_clk(i_clk));
Mul0000000001  u_0000000123_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[24*12+:12]), .o_data(C[24][0]), .i_clk(i_clk));
Mul0000000001  u_0000000124_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[280*12+:12]), .o_data(A[24][1]), .i_clk(i_clk));
Mul0000000001  u_0000000125_Mul0000000001(.i_data_1(c_plus_d[24][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[24][1]), .i_clk(i_clk));
Mul0000000001  u_0000000126_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[280*12+:12]), .o_data(C[24][1]), .i_clk(i_clk));
Mul0000000001  u_0000000127_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[536*12+:12]), .o_data(A[24][2]), .i_clk(i_clk));
Mul0000000001  u_0000000128_Mul0000000001(.i_data_1(c_plus_d[24][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[24][2]), .i_clk(i_clk));
Mul0000000001  u_0000000129_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[536*12+:12]), .o_data(C[24][2]), .i_clk(i_clk));
Mul0000000001  u_000000012A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[792*12+:12]), .o_data(A[24][3]), .i_clk(i_clk));
Mul0000000001  u_000000012B_Mul0000000001(.i_data_1(c_plus_d[24][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[24][3]), .i_clk(i_clk));
Mul0000000001  u_000000012C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[792*12+:12]), .o_data(C[24][3]), .i_clk(i_clk));
Mul0000000001  u_000000012D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[25*12+:12]), .o_data(A[25][0]), .i_clk(i_clk));
Mul0000000001  u_000000012E_Mul0000000001(.i_data_1(c_plus_d[25][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[25][0]), .i_clk(i_clk));
Mul0000000001  u_000000012F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[25*12+:12]), .o_data(C[25][0]), .i_clk(i_clk));
Mul0000000001  u_0000000130_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[281*12+:12]), .o_data(A[25][1]), .i_clk(i_clk));
Mul0000000001  u_0000000131_Mul0000000001(.i_data_1(c_plus_d[25][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[25][1]), .i_clk(i_clk));
Mul0000000001  u_0000000132_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[281*12+:12]), .o_data(C[25][1]), .i_clk(i_clk));
Mul0000000001  u_0000000133_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[537*12+:12]), .o_data(A[25][2]), .i_clk(i_clk));
Mul0000000001  u_0000000134_Mul0000000001(.i_data_1(c_plus_d[25][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[25][2]), .i_clk(i_clk));
Mul0000000001  u_0000000135_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[537*12+:12]), .o_data(C[25][2]), .i_clk(i_clk));
Mul0000000001  u_0000000136_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[793*12+:12]), .o_data(A[25][3]), .i_clk(i_clk));
Mul0000000001  u_0000000137_Mul0000000001(.i_data_1(c_plus_d[25][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[25][3]), .i_clk(i_clk));
Mul0000000001  u_0000000138_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[793*12+:12]), .o_data(C[25][3]), .i_clk(i_clk));
Mul0000000001  u_0000000139_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[26*12+:12]), .o_data(A[26][0]), .i_clk(i_clk));
Mul0000000001  u_000000013A_Mul0000000001(.i_data_1(c_plus_d[26][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[26][0]), .i_clk(i_clk));
Mul0000000001  u_000000013B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[26*12+:12]), .o_data(C[26][0]), .i_clk(i_clk));
Mul0000000001  u_000000013C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[282*12+:12]), .o_data(A[26][1]), .i_clk(i_clk));
Mul0000000001  u_000000013D_Mul0000000001(.i_data_1(c_plus_d[26][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[26][1]), .i_clk(i_clk));
Mul0000000001  u_000000013E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[282*12+:12]), .o_data(C[26][1]), .i_clk(i_clk));
Mul0000000001  u_000000013F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[538*12+:12]), .o_data(A[26][2]), .i_clk(i_clk));
Mul0000000001  u_0000000140_Mul0000000001(.i_data_1(c_plus_d[26][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[26][2]), .i_clk(i_clk));
Mul0000000001  u_0000000141_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[538*12+:12]), .o_data(C[26][2]), .i_clk(i_clk));
Mul0000000001  u_0000000142_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[794*12+:12]), .o_data(A[26][3]), .i_clk(i_clk));
Mul0000000001  u_0000000143_Mul0000000001(.i_data_1(c_plus_d[26][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[26][3]), .i_clk(i_clk));
Mul0000000001  u_0000000144_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[794*12+:12]), .o_data(C[26][3]), .i_clk(i_clk));
Mul0000000001  u_0000000145_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[27*12+:12]), .o_data(A[27][0]), .i_clk(i_clk));
Mul0000000001  u_0000000146_Mul0000000001(.i_data_1(c_plus_d[27][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[27][0]), .i_clk(i_clk));
Mul0000000001  u_0000000147_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[27*12+:12]), .o_data(C[27][0]), .i_clk(i_clk));
Mul0000000001  u_0000000148_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[283*12+:12]), .o_data(A[27][1]), .i_clk(i_clk));
Mul0000000001  u_0000000149_Mul0000000001(.i_data_1(c_plus_d[27][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[27][1]), .i_clk(i_clk));
Mul0000000001  u_000000014A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[283*12+:12]), .o_data(C[27][1]), .i_clk(i_clk));
Mul0000000001  u_000000014B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[539*12+:12]), .o_data(A[27][2]), .i_clk(i_clk));
Mul0000000001  u_000000014C_Mul0000000001(.i_data_1(c_plus_d[27][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[27][2]), .i_clk(i_clk));
Mul0000000001  u_000000014D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[539*12+:12]), .o_data(C[27][2]), .i_clk(i_clk));
Mul0000000001  u_000000014E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[795*12+:12]), .o_data(A[27][3]), .i_clk(i_clk));
Mul0000000001  u_000000014F_Mul0000000001(.i_data_1(c_plus_d[27][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[27][3]), .i_clk(i_clk));
Mul0000000001  u_0000000150_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[795*12+:12]), .o_data(C[27][3]), .i_clk(i_clk));
Mul0000000001  u_0000000151_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[28*12+:12]), .o_data(A[28][0]), .i_clk(i_clk));
Mul0000000001  u_0000000152_Mul0000000001(.i_data_1(c_plus_d[28][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[28][0]), .i_clk(i_clk));
Mul0000000001  u_0000000153_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[28*12+:12]), .o_data(C[28][0]), .i_clk(i_clk));
Mul0000000001  u_0000000154_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[284*12+:12]), .o_data(A[28][1]), .i_clk(i_clk));
Mul0000000001  u_0000000155_Mul0000000001(.i_data_1(c_plus_d[28][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[28][1]), .i_clk(i_clk));
Mul0000000001  u_0000000156_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[284*12+:12]), .o_data(C[28][1]), .i_clk(i_clk));
Mul0000000001  u_0000000157_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[540*12+:12]), .o_data(A[28][2]), .i_clk(i_clk));
Mul0000000001  u_0000000158_Mul0000000001(.i_data_1(c_plus_d[28][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[28][2]), .i_clk(i_clk));
Mul0000000001  u_0000000159_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[540*12+:12]), .o_data(C[28][2]), .i_clk(i_clk));
Mul0000000001  u_000000015A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[796*12+:12]), .o_data(A[28][3]), .i_clk(i_clk));
Mul0000000001  u_000000015B_Mul0000000001(.i_data_1(c_plus_d[28][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[28][3]), .i_clk(i_clk));
Mul0000000001  u_000000015C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[796*12+:12]), .o_data(C[28][3]), .i_clk(i_clk));
Mul0000000001  u_000000015D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[29*12+:12]), .o_data(A[29][0]), .i_clk(i_clk));
Mul0000000001  u_000000015E_Mul0000000001(.i_data_1(c_plus_d[29][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[29][0]), .i_clk(i_clk));
Mul0000000001  u_000000015F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[29*12+:12]), .o_data(C[29][0]), .i_clk(i_clk));
Mul0000000001  u_0000000160_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[285*12+:12]), .o_data(A[29][1]), .i_clk(i_clk));
Mul0000000001  u_0000000161_Mul0000000001(.i_data_1(c_plus_d[29][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[29][1]), .i_clk(i_clk));
Mul0000000001  u_0000000162_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[285*12+:12]), .o_data(C[29][1]), .i_clk(i_clk));
Mul0000000001  u_0000000163_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[541*12+:12]), .o_data(A[29][2]), .i_clk(i_clk));
Mul0000000001  u_0000000164_Mul0000000001(.i_data_1(c_plus_d[29][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[29][2]), .i_clk(i_clk));
Mul0000000001  u_0000000165_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[541*12+:12]), .o_data(C[29][2]), .i_clk(i_clk));
Mul0000000001  u_0000000166_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[797*12+:12]), .o_data(A[29][3]), .i_clk(i_clk));
Mul0000000001  u_0000000167_Mul0000000001(.i_data_1(c_plus_d[29][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[29][3]), .i_clk(i_clk));
Mul0000000001  u_0000000168_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[797*12+:12]), .o_data(C[29][3]), .i_clk(i_clk));
Mul0000000001  u_0000000169_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[30*12+:12]), .o_data(A[30][0]), .i_clk(i_clk));
Mul0000000001  u_000000016A_Mul0000000001(.i_data_1(c_plus_d[30][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[30][0]), .i_clk(i_clk));
Mul0000000001  u_000000016B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[30*12+:12]), .o_data(C[30][0]), .i_clk(i_clk));
Mul0000000001  u_000000016C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[286*12+:12]), .o_data(A[30][1]), .i_clk(i_clk));
Mul0000000001  u_000000016D_Mul0000000001(.i_data_1(c_plus_d[30][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[30][1]), .i_clk(i_clk));
Mul0000000001  u_000000016E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[286*12+:12]), .o_data(C[30][1]), .i_clk(i_clk));
Mul0000000001  u_000000016F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[542*12+:12]), .o_data(A[30][2]), .i_clk(i_clk));
Mul0000000001  u_0000000170_Mul0000000001(.i_data_1(c_plus_d[30][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[30][2]), .i_clk(i_clk));
Mul0000000001  u_0000000171_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[542*12+:12]), .o_data(C[30][2]), .i_clk(i_clk));
Mul0000000001  u_0000000172_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[798*12+:12]), .o_data(A[30][3]), .i_clk(i_clk));
Mul0000000001  u_0000000173_Mul0000000001(.i_data_1(c_plus_d[30][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[30][3]), .i_clk(i_clk));
Mul0000000001  u_0000000174_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[798*12+:12]), .o_data(C[30][3]), .i_clk(i_clk));
Mul0000000001  u_0000000175_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[31*12+:12]), .o_data(A[31][0]), .i_clk(i_clk));
Mul0000000001  u_0000000176_Mul0000000001(.i_data_1(c_plus_d[31][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[31][0]), .i_clk(i_clk));
Mul0000000001  u_0000000177_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[31*12+:12]), .o_data(C[31][0]), .i_clk(i_clk));
Mul0000000001  u_0000000178_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[287*12+:12]), .o_data(A[31][1]), .i_clk(i_clk));
Mul0000000001  u_0000000179_Mul0000000001(.i_data_1(c_plus_d[31][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[31][1]), .i_clk(i_clk));
Mul0000000001  u_000000017A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[287*12+:12]), .o_data(C[31][1]), .i_clk(i_clk));
Mul0000000001  u_000000017B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[543*12+:12]), .o_data(A[31][2]), .i_clk(i_clk));
Mul0000000001  u_000000017C_Mul0000000001(.i_data_1(c_plus_d[31][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[31][2]), .i_clk(i_clk));
Mul0000000001  u_000000017D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[543*12+:12]), .o_data(C[31][2]), .i_clk(i_clk));
Mul0000000001  u_000000017E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[799*12+:12]), .o_data(A[31][3]), .i_clk(i_clk));
Mul0000000001  u_000000017F_Mul0000000001(.i_data_1(c_plus_d[31][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[31][3]), .i_clk(i_clk));
Mul0000000001  u_0000000180_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[799*12+:12]), .o_data(C[31][3]), .i_clk(i_clk));
Mul0000000001  u_0000000181_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[32*12+:12]), .o_data(A[32][0]), .i_clk(i_clk));
Mul0000000001  u_0000000182_Mul0000000001(.i_data_1(c_plus_d[32][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[32][0]), .i_clk(i_clk));
Mul0000000001  u_0000000183_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[32*12+:12]), .o_data(C[32][0]), .i_clk(i_clk));
Mul0000000001  u_0000000184_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[288*12+:12]), .o_data(A[32][1]), .i_clk(i_clk));
Mul0000000001  u_0000000185_Mul0000000001(.i_data_1(c_plus_d[32][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[32][1]), .i_clk(i_clk));
Mul0000000001  u_0000000186_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[288*12+:12]), .o_data(C[32][1]), .i_clk(i_clk));
Mul0000000001  u_0000000187_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[544*12+:12]), .o_data(A[32][2]), .i_clk(i_clk));
Mul0000000001  u_0000000188_Mul0000000001(.i_data_1(c_plus_d[32][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[32][2]), .i_clk(i_clk));
Mul0000000001  u_0000000189_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[544*12+:12]), .o_data(C[32][2]), .i_clk(i_clk));
Mul0000000001  u_000000018A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[800*12+:12]), .o_data(A[32][3]), .i_clk(i_clk));
Mul0000000001  u_000000018B_Mul0000000001(.i_data_1(c_plus_d[32][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[32][3]), .i_clk(i_clk));
Mul0000000001  u_000000018C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[800*12+:12]), .o_data(C[32][3]), .i_clk(i_clk));
Mul0000000001  u_000000018D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[33*12+:12]), .o_data(A[33][0]), .i_clk(i_clk));
Mul0000000001  u_000000018E_Mul0000000001(.i_data_1(c_plus_d[33][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[33][0]), .i_clk(i_clk));
Mul0000000001  u_000000018F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[33*12+:12]), .o_data(C[33][0]), .i_clk(i_clk));
Mul0000000001  u_0000000190_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[289*12+:12]), .o_data(A[33][1]), .i_clk(i_clk));
Mul0000000001  u_0000000191_Mul0000000001(.i_data_1(c_plus_d[33][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[33][1]), .i_clk(i_clk));
Mul0000000001  u_0000000192_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[289*12+:12]), .o_data(C[33][1]), .i_clk(i_clk));
Mul0000000001  u_0000000193_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[545*12+:12]), .o_data(A[33][2]), .i_clk(i_clk));
Mul0000000001  u_0000000194_Mul0000000001(.i_data_1(c_plus_d[33][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[33][2]), .i_clk(i_clk));
Mul0000000001  u_0000000195_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[545*12+:12]), .o_data(C[33][2]), .i_clk(i_clk));
Mul0000000001  u_0000000196_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[801*12+:12]), .o_data(A[33][3]), .i_clk(i_clk));
Mul0000000001  u_0000000197_Mul0000000001(.i_data_1(c_plus_d[33][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[33][3]), .i_clk(i_clk));
Mul0000000001  u_0000000198_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[801*12+:12]), .o_data(C[33][3]), .i_clk(i_clk));
Mul0000000001  u_0000000199_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[34*12+:12]), .o_data(A[34][0]), .i_clk(i_clk));
Mul0000000001  u_000000019A_Mul0000000001(.i_data_1(c_plus_d[34][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[34][0]), .i_clk(i_clk));
Mul0000000001  u_000000019B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[34*12+:12]), .o_data(C[34][0]), .i_clk(i_clk));
Mul0000000001  u_000000019C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[290*12+:12]), .o_data(A[34][1]), .i_clk(i_clk));
Mul0000000001  u_000000019D_Mul0000000001(.i_data_1(c_plus_d[34][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[34][1]), .i_clk(i_clk));
Mul0000000001  u_000000019E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[290*12+:12]), .o_data(C[34][1]), .i_clk(i_clk));
Mul0000000001  u_000000019F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[546*12+:12]), .o_data(A[34][2]), .i_clk(i_clk));
Mul0000000001  u_00000001A0_Mul0000000001(.i_data_1(c_plus_d[34][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[34][2]), .i_clk(i_clk));
Mul0000000001  u_00000001A1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[546*12+:12]), .o_data(C[34][2]), .i_clk(i_clk));
Mul0000000001  u_00000001A2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[802*12+:12]), .o_data(A[34][3]), .i_clk(i_clk));
Mul0000000001  u_00000001A3_Mul0000000001(.i_data_1(c_plus_d[34][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[34][3]), .i_clk(i_clk));
Mul0000000001  u_00000001A4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[802*12+:12]), .o_data(C[34][3]), .i_clk(i_clk));
Mul0000000001  u_00000001A5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[35*12+:12]), .o_data(A[35][0]), .i_clk(i_clk));
Mul0000000001  u_00000001A6_Mul0000000001(.i_data_1(c_plus_d[35][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[35][0]), .i_clk(i_clk));
Mul0000000001  u_00000001A7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[35*12+:12]), .o_data(C[35][0]), .i_clk(i_clk));
Mul0000000001  u_00000001A8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[291*12+:12]), .o_data(A[35][1]), .i_clk(i_clk));
Mul0000000001  u_00000001A9_Mul0000000001(.i_data_1(c_plus_d[35][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[35][1]), .i_clk(i_clk));
Mul0000000001  u_00000001AA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[291*12+:12]), .o_data(C[35][1]), .i_clk(i_clk));
Mul0000000001  u_00000001AB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[547*12+:12]), .o_data(A[35][2]), .i_clk(i_clk));
Mul0000000001  u_00000001AC_Mul0000000001(.i_data_1(c_plus_d[35][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[35][2]), .i_clk(i_clk));
Mul0000000001  u_00000001AD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[547*12+:12]), .o_data(C[35][2]), .i_clk(i_clk));
Mul0000000001  u_00000001AE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[803*12+:12]), .o_data(A[35][3]), .i_clk(i_clk));
Mul0000000001  u_00000001AF_Mul0000000001(.i_data_1(c_plus_d[35][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[35][3]), .i_clk(i_clk));
Mul0000000001  u_00000001B0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[803*12+:12]), .o_data(C[35][3]), .i_clk(i_clk));
Mul0000000001  u_00000001B1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[36*12+:12]), .o_data(A[36][0]), .i_clk(i_clk));
Mul0000000001  u_00000001B2_Mul0000000001(.i_data_1(c_plus_d[36][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[36][0]), .i_clk(i_clk));
Mul0000000001  u_00000001B3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[36*12+:12]), .o_data(C[36][0]), .i_clk(i_clk));
Mul0000000001  u_00000001B4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[292*12+:12]), .o_data(A[36][1]), .i_clk(i_clk));
Mul0000000001  u_00000001B5_Mul0000000001(.i_data_1(c_plus_d[36][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[36][1]), .i_clk(i_clk));
Mul0000000001  u_00000001B6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[292*12+:12]), .o_data(C[36][1]), .i_clk(i_clk));
Mul0000000001  u_00000001B7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[548*12+:12]), .o_data(A[36][2]), .i_clk(i_clk));
Mul0000000001  u_00000001B8_Mul0000000001(.i_data_1(c_plus_d[36][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[36][2]), .i_clk(i_clk));
Mul0000000001  u_00000001B9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[548*12+:12]), .o_data(C[36][2]), .i_clk(i_clk));
Mul0000000001  u_00000001BA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[804*12+:12]), .o_data(A[36][3]), .i_clk(i_clk));
Mul0000000001  u_00000001BB_Mul0000000001(.i_data_1(c_plus_d[36][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[36][3]), .i_clk(i_clk));
Mul0000000001  u_00000001BC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[804*12+:12]), .o_data(C[36][3]), .i_clk(i_clk));
Mul0000000001  u_00000001BD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[37*12+:12]), .o_data(A[37][0]), .i_clk(i_clk));
Mul0000000001  u_00000001BE_Mul0000000001(.i_data_1(c_plus_d[37][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[37][0]), .i_clk(i_clk));
Mul0000000001  u_00000001BF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[37*12+:12]), .o_data(C[37][0]), .i_clk(i_clk));
Mul0000000001  u_00000001C0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[293*12+:12]), .o_data(A[37][1]), .i_clk(i_clk));
Mul0000000001  u_00000001C1_Mul0000000001(.i_data_1(c_plus_d[37][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[37][1]), .i_clk(i_clk));
Mul0000000001  u_00000001C2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[293*12+:12]), .o_data(C[37][1]), .i_clk(i_clk));
Mul0000000001  u_00000001C3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[549*12+:12]), .o_data(A[37][2]), .i_clk(i_clk));
Mul0000000001  u_00000001C4_Mul0000000001(.i_data_1(c_plus_d[37][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[37][2]), .i_clk(i_clk));
Mul0000000001  u_00000001C5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[549*12+:12]), .o_data(C[37][2]), .i_clk(i_clk));
Mul0000000001  u_00000001C6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[805*12+:12]), .o_data(A[37][3]), .i_clk(i_clk));
Mul0000000001  u_00000001C7_Mul0000000001(.i_data_1(c_plus_d[37][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[37][3]), .i_clk(i_clk));
Mul0000000001  u_00000001C8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[805*12+:12]), .o_data(C[37][3]), .i_clk(i_clk));
Mul0000000001  u_00000001C9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[38*12+:12]), .o_data(A[38][0]), .i_clk(i_clk));
Mul0000000001  u_00000001CA_Mul0000000001(.i_data_1(c_plus_d[38][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[38][0]), .i_clk(i_clk));
Mul0000000001  u_00000001CB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[38*12+:12]), .o_data(C[38][0]), .i_clk(i_clk));
Mul0000000001  u_00000001CC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[294*12+:12]), .o_data(A[38][1]), .i_clk(i_clk));
Mul0000000001  u_00000001CD_Mul0000000001(.i_data_1(c_plus_d[38][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[38][1]), .i_clk(i_clk));
Mul0000000001  u_00000001CE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[294*12+:12]), .o_data(C[38][1]), .i_clk(i_clk));
Mul0000000001  u_00000001CF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[550*12+:12]), .o_data(A[38][2]), .i_clk(i_clk));
Mul0000000001  u_00000001D0_Mul0000000001(.i_data_1(c_plus_d[38][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[38][2]), .i_clk(i_clk));
Mul0000000001  u_00000001D1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[550*12+:12]), .o_data(C[38][2]), .i_clk(i_clk));
Mul0000000001  u_00000001D2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[806*12+:12]), .o_data(A[38][3]), .i_clk(i_clk));
Mul0000000001  u_00000001D3_Mul0000000001(.i_data_1(c_plus_d[38][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[38][3]), .i_clk(i_clk));
Mul0000000001  u_00000001D4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[806*12+:12]), .o_data(C[38][3]), .i_clk(i_clk));
Mul0000000001  u_00000001D5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[39*12+:12]), .o_data(A[39][0]), .i_clk(i_clk));
Mul0000000001  u_00000001D6_Mul0000000001(.i_data_1(c_plus_d[39][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[39][0]), .i_clk(i_clk));
Mul0000000001  u_00000001D7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[39*12+:12]), .o_data(C[39][0]), .i_clk(i_clk));
Mul0000000001  u_00000001D8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[295*12+:12]), .o_data(A[39][1]), .i_clk(i_clk));
Mul0000000001  u_00000001D9_Mul0000000001(.i_data_1(c_plus_d[39][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[39][1]), .i_clk(i_clk));
Mul0000000001  u_00000001DA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[295*12+:12]), .o_data(C[39][1]), .i_clk(i_clk));
Mul0000000001  u_00000001DB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[551*12+:12]), .o_data(A[39][2]), .i_clk(i_clk));
Mul0000000001  u_00000001DC_Mul0000000001(.i_data_1(c_plus_d[39][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[39][2]), .i_clk(i_clk));
Mul0000000001  u_00000001DD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[551*12+:12]), .o_data(C[39][2]), .i_clk(i_clk));
Mul0000000001  u_00000001DE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[807*12+:12]), .o_data(A[39][3]), .i_clk(i_clk));
Mul0000000001  u_00000001DF_Mul0000000001(.i_data_1(c_plus_d[39][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[39][3]), .i_clk(i_clk));
Mul0000000001  u_00000001E0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[807*12+:12]), .o_data(C[39][3]), .i_clk(i_clk));
Mul0000000001  u_00000001E1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[40*12+:12]), .o_data(A[40][0]), .i_clk(i_clk));
Mul0000000001  u_00000001E2_Mul0000000001(.i_data_1(c_plus_d[40][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[40][0]), .i_clk(i_clk));
Mul0000000001  u_00000001E3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[40*12+:12]), .o_data(C[40][0]), .i_clk(i_clk));
Mul0000000001  u_00000001E4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[296*12+:12]), .o_data(A[40][1]), .i_clk(i_clk));
Mul0000000001  u_00000001E5_Mul0000000001(.i_data_1(c_plus_d[40][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[40][1]), .i_clk(i_clk));
Mul0000000001  u_00000001E6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[296*12+:12]), .o_data(C[40][1]), .i_clk(i_clk));
Mul0000000001  u_00000001E7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[552*12+:12]), .o_data(A[40][2]), .i_clk(i_clk));
Mul0000000001  u_00000001E8_Mul0000000001(.i_data_1(c_plus_d[40][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[40][2]), .i_clk(i_clk));
Mul0000000001  u_00000001E9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[552*12+:12]), .o_data(C[40][2]), .i_clk(i_clk));
Mul0000000001  u_00000001EA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[808*12+:12]), .o_data(A[40][3]), .i_clk(i_clk));
Mul0000000001  u_00000001EB_Mul0000000001(.i_data_1(c_plus_d[40][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[40][3]), .i_clk(i_clk));
Mul0000000001  u_00000001EC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[808*12+:12]), .o_data(C[40][3]), .i_clk(i_clk));
Mul0000000001  u_00000001ED_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[41*12+:12]), .o_data(A[41][0]), .i_clk(i_clk));
Mul0000000001  u_00000001EE_Mul0000000001(.i_data_1(c_plus_d[41][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[41][0]), .i_clk(i_clk));
Mul0000000001  u_00000001EF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[41*12+:12]), .o_data(C[41][0]), .i_clk(i_clk));
Mul0000000001  u_00000001F0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[297*12+:12]), .o_data(A[41][1]), .i_clk(i_clk));
Mul0000000001  u_00000001F1_Mul0000000001(.i_data_1(c_plus_d[41][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[41][1]), .i_clk(i_clk));
Mul0000000001  u_00000001F2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[297*12+:12]), .o_data(C[41][1]), .i_clk(i_clk));
Mul0000000001  u_00000001F3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[553*12+:12]), .o_data(A[41][2]), .i_clk(i_clk));
Mul0000000001  u_00000001F4_Mul0000000001(.i_data_1(c_plus_d[41][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[41][2]), .i_clk(i_clk));
Mul0000000001  u_00000001F5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[553*12+:12]), .o_data(C[41][2]), .i_clk(i_clk));
Mul0000000001  u_00000001F6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[809*12+:12]), .o_data(A[41][3]), .i_clk(i_clk));
Mul0000000001  u_00000001F7_Mul0000000001(.i_data_1(c_plus_d[41][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[41][3]), .i_clk(i_clk));
Mul0000000001  u_00000001F8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[809*12+:12]), .o_data(C[41][3]), .i_clk(i_clk));
Mul0000000001  u_00000001F9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[42*12+:12]), .o_data(A[42][0]), .i_clk(i_clk));
Mul0000000001  u_00000001FA_Mul0000000001(.i_data_1(c_plus_d[42][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[42][0]), .i_clk(i_clk));
Mul0000000001  u_00000001FB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[42*12+:12]), .o_data(C[42][0]), .i_clk(i_clk));
Mul0000000001  u_00000001FC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[298*12+:12]), .o_data(A[42][1]), .i_clk(i_clk));
Mul0000000001  u_00000001FD_Mul0000000001(.i_data_1(c_plus_d[42][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[42][1]), .i_clk(i_clk));
Mul0000000001  u_00000001FE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[298*12+:12]), .o_data(C[42][1]), .i_clk(i_clk));
Mul0000000001  u_00000001FF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[554*12+:12]), .o_data(A[42][2]), .i_clk(i_clk));
Mul0000000001  u_0000000200_Mul0000000001(.i_data_1(c_plus_d[42][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[42][2]), .i_clk(i_clk));
Mul0000000001  u_0000000201_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[554*12+:12]), .o_data(C[42][2]), .i_clk(i_clk));
Mul0000000001  u_0000000202_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[810*12+:12]), .o_data(A[42][3]), .i_clk(i_clk));
Mul0000000001  u_0000000203_Mul0000000001(.i_data_1(c_plus_d[42][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[42][3]), .i_clk(i_clk));
Mul0000000001  u_0000000204_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[810*12+:12]), .o_data(C[42][3]), .i_clk(i_clk));
Mul0000000001  u_0000000205_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[43*12+:12]), .o_data(A[43][0]), .i_clk(i_clk));
Mul0000000001  u_0000000206_Mul0000000001(.i_data_1(c_plus_d[43][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[43][0]), .i_clk(i_clk));
Mul0000000001  u_0000000207_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[43*12+:12]), .o_data(C[43][0]), .i_clk(i_clk));
Mul0000000001  u_0000000208_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[299*12+:12]), .o_data(A[43][1]), .i_clk(i_clk));
Mul0000000001  u_0000000209_Mul0000000001(.i_data_1(c_plus_d[43][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[43][1]), .i_clk(i_clk));
Mul0000000001  u_000000020A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[299*12+:12]), .o_data(C[43][1]), .i_clk(i_clk));
Mul0000000001  u_000000020B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[555*12+:12]), .o_data(A[43][2]), .i_clk(i_clk));
Mul0000000001  u_000000020C_Mul0000000001(.i_data_1(c_plus_d[43][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[43][2]), .i_clk(i_clk));
Mul0000000001  u_000000020D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[555*12+:12]), .o_data(C[43][2]), .i_clk(i_clk));
Mul0000000001  u_000000020E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[811*12+:12]), .o_data(A[43][3]), .i_clk(i_clk));
Mul0000000001  u_000000020F_Mul0000000001(.i_data_1(c_plus_d[43][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[43][3]), .i_clk(i_clk));
Mul0000000001  u_0000000210_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[811*12+:12]), .o_data(C[43][3]), .i_clk(i_clk));
Mul0000000001  u_0000000211_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[44*12+:12]), .o_data(A[44][0]), .i_clk(i_clk));
Mul0000000001  u_0000000212_Mul0000000001(.i_data_1(c_plus_d[44][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[44][0]), .i_clk(i_clk));
Mul0000000001  u_0000000213_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[44*12+:12]), .o_data(C[44][0]), .i_clk(i_clk));
Mul0000000001  u_0000000214_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[300*12+:12]), .o_data(A[44][1]), .i_clk(i_clk));
Mul0000000001  u_0000000215_Mul0000000001(.i_data_1(c_plus_d[44][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[44][1]), .i_clk(i_clk));
Mul0000000001  u_0000000216_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[300*12+:12]), .o_data(C[44][1]), .i_clk(i_clk));
Mul0000000001  u_0000000217_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[556*12+:12]), .o_data(A[44][2]), .i_clk(i_clk));
Mul0000000001  u_0000000218_Mul0000000001(.i_data_1(c_plus_d[44][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[44][2]), .i_clk(i_clk));
Mul0000000001  u_0000000219_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[556*12+:12]), .o_data(C[44][2]), .i_clk(i_clk));
Mul0000000001  u_000000021A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[812*12+:12]), .o_data(A[44][3]), .i_clk(i_clk));
Mul0000000001  u_000000021B_Mul0000000001(.i_data_1(c_plus_d[44][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[44][3]), .i_clk(i_clk));
Mul0000000001  u_000000021C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[812*12+:12]), .o_data(C[44][3]), .i_clk(i_clk));
Mul0000000001  u_000000021D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[45*12+:12]), .o_data(A[45][0]), .i_clk(i_clk));
Mul0000000001  u_000000021E_Mul0000000001(.i_data_1(c_plus_d[45][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[45][0]), .i_clk(i_clk));
Mul0000000001  u_000000021F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[45*12+:12]), .o_data(C[45][0]), .i_clk(i_clk));
Mul0000000001  u_0000000220_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[301*12+:12]), .o_data(A[45][1]), .i_clk(i_clk));
Mul0000000001  u_0000000221_Mul0000000001(.i_data_1(c_plus_d[45][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[45][1]), .i_clk(i_clk));
Mul0000000001  u_0000000222_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[301*12+:12]), .o_data(C[45][1]), .i_clk(i_clk));
Mul0000000001  u_0000000223_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[557*12+:12]), .o_data(A[45][2]), .i_clk(i_clk));
Mul0000000001  u_0000000224_Mul0000000001(.i_data_1(c_plus_d[45][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[45][2]), .i_clk(i_clk));
Mul0000000001  u_0000000225_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[557*12+:12]), .o_data(C[45][2]), .i_clk(i_clk));
Mul0000000001  u_0000000226_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[813*12+:12]), .o_data(A[45][3]), .i_clk(i_clk));
Mul0000000001  u_0000000227_Mul0000000001(.i_data_1(c_plus_d[45][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[45][3]), .i_clk(i_clk));
Mul0000000001  u_0000000228_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[813*12+:12]), .o_data(C[45][3]), .i_clk(i_clk));
Mul0000000001  u_0000000229_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[46*12+:12]), .o_data(A[46][0]), .i_clk(i_clk));
Mul0000000001  u_000000022A_Mul0000000001(.i_data_1(c_plus_d[46][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[46][0]), .i_clk(i_clk));
Mul0000000001  u_000000022B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[46*12+:12]), .o_data(C[46][0]), .i_clk(i_clk));
Mul0000000001  u_000000022C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[302*12+:12]), .o_data(A[46][1]), .i_clk(i_clk));
Mul0000000001  u_000000022D_Mul0000000001(.i_data_1(c_plus_d[46][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[46][1]), .i_clk(i_clk));
Mul0000000001  u_000000022E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[302*12+:12]), .o_data(C[46][1]), .i_clk(i_clk));
Mul0000000001  u_000000022F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[558*12+:12]), .o_data(A[46][2]), .i_clk(i_clk));
Mul0000000001  u_0000000230_Mul0000000001(.i_data_1(c_plus_d[46][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[46][2]), .i_clk(i_clk));
Mul0000000001  u_0000000231_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[558*12+:12]), .o_data(C[46][2]), .i_clk(i_clk));
Mul0000000001  u_0000000232_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[814*12+:12]), .o_data(A[46][3]), .i_clk(i_clk));
Mul0000000001  u_0000000233_Mul0000000001(.i_data_1(c_plus_d[46][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[46][3]), .i_clk(i_clk));
Mul0000000001  u_0000000234_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[814*12+:12]), .o_data(C[46][3]), .i_clk(i_clk));
Mul0000000001  u_0000000235_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[47*12+:12]), .o_data(A[47][0]), .i_clk(i_clk));
Mul0000000001  u_0000000236_Mul0000000001(.i_data_1(c_plus_d[47][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[47][0]), .i_clk(i_clk));
Mul0000000001  u_0000000237_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[47*12+:12]), .o_data(C[47][0]), .i_clk(i_clk));
Mul0000000001  u_0000000238_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[303*12+:12]), .o_data(A[47][1]), .i_clk(i_clk));
Mul0000000001  u_0000000239_Mul0000000001(.i_data_1(c_plus_d[47][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[47][1]), .i_clk(i_clk));
Mul0000000001  u_000000023A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[303*12+:12]), .o_data(C[47][1]), .i_clk(i_clk));
Mul0000000001  u_000000023B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[559*12+:12]), .o_data(A[47][2]), .i_clk(i_clk));
Mul0000000001  u_000000023C_Mul0000000001(.i_data_1(c_plus_d[47][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[47][2]), .i_clk(i_clk));
Mul0000000001  u_000000023D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[559*12+:12]), .o_data(C[47][2]), .i_clk(i_clk));
Mul0000000001  u_000000023E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[815*12+:12]), .o_data(A[47][3]), .i_clk(i_clk));
Mul0000000001  u_000000023F_Mul0000000001(.i_data_1(c_plus_d[47][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[47][3]), .i_clk(i_clk));
Mul0000000001  u_0000000240_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[815*12+:12]), .o_data(C[47][3]), .i_clk(i_clk));
Mul0000000001  u_0000000241_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[48*12+:12]), .o_data(A[48][0]), .i_clk(i_clk));
Mul0000000001  u_0000000242_Mul0000000001(.i_data_1(c_plus_d[48][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[48][0]), .i_clk(i_clk));
Mul0000000001  u_0000000243_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[48*12+:12]), .o_data(C[48][0]), .i_clk(i_clk));
Mul0000000001  u_0000000244_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[304*12+:12]), .o_data(A[48][1]), .i_clk(i_clk));
Mul0000000001  u_0000000245_Mul0000000001(.i_data_1(c_plus_d[48][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[48][1]), .i_clk(i_clk));
Mul0000000001  u_0000000246_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[304*12+:12]), .o_data(C[48][1]), .i_clk(i_clk));
Mul0000000001  u_0000000247_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[560*12+:12]), .o_data(A[48][2]), .i_clk(i_clk));
Mul0000000001  u_0000000248_Mul0000000001(.i_data_1(c_plus_d[48][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[48][2]), .i_clk(i_clk));
Mul0000000001  u_0000000249_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[560*12+:12]), .o_data(C[48][2]), .i_clk(i_clk));
Mul0000000001  u_000000024A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[816*12+:12]), .o_data(A[48][3]), .i_clk(i_clk));
Mul0000000001  u_000000024B_Mul0000000001(.i_data_1(c_plus_d[48][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[48][3]), .i_clk(i_clk));
Mul0000000001  u_000000024C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[816*12+:12]), .o_data(C[48][3]), .i_clk(i_clk));
Mul0000000001  u_000000024D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[49*12+:12]), .o_data(A[49][0]), .i_clk(i_clk));
Mul0000000001  u_000000024E_Mul0000000001(.i_data_1(c_plus_d[49][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[49][0]), .i_clk(i_clk));
Mul0000000001  u_000000024F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[49*12+:12]), .o_data(C[49][0]), .i_clk(i_clk));
Mul0000000001  u_0000000250_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[305*12+:12]), .o_data(A[49][1]), .i_clk(i_clk));
Mul0000000001  u_0000000251_Mul0000000001(.i_data_1(c_plus_d[49][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[49][1]), .i_clk(i_clk));
Mul0000000001  u_0000000252_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[305*12+:12]), .o_data(C[49][1]), .i_clk(i_clk));
Mul0000000001  u_0000000253_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[561*12+:12]), .o_data(A[49][2]), .i_clk(i_clk));
Mul0000000001  u_0000000254_Mul0000000001(.i_data_1(c_plus_d[49][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[49][2]), .i_clk(i_clk));
Mul0000000001  u_0000000255_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[561*12+:12]), .o_data(C[49][2]), .i_clk(i_clk));
Mul0000000001  u_0000000256_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[817*12+:12]), .o_data(A[49][3]), .i_clk(i_clk));
Mul0000000001  u_0000000257_Mul0000000001(.i_data_1(c_plus_d[49][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[49][3]), .i_clk(i_clk));
Mul0000000001  u_0000000258_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[817*12+:12]), .o_data(C[49][3]), .i_clk(i_clk));
Mul0000000001  u_0000000259_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[50*12+:12]), .o_data(A[50][0]), .i_clk(i_clk));
Mul0000000001  u_000000025A_Mul0000000001(.i_data_1(c_plus_d[50][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[50][0]), .i_clk(i_clk));
Mul0000000001  u_000000025B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[50*12+:12]), .o_data(C[50][0]), .i_clk(i_clk));
Mul0000000001  u_000000025C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[306*12+:12]), .o_data(A[50][1]), .i_clk(i_clk));
Mul0000000001  u_000000025D_Mul0000000001(.i_data_1(c_plus_d[50][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[50][1]), .i_clk(i_clk));
Mul0000000001  u_000000025E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[306*12+:12]), .o_data(C[50][1]), .i_clk(i_clk));
Mul0000000001  u_000000025F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[562*12+:12]), .o_data(A[50][2]), .i_clk(i_clk));
Mul0000000001  u_0000000260_Mul0000000001(.i_data_1(c_plus_d[50][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[50][2]), .i_clk(i_clk));
Mul0000000001  u_0000000261_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[562*12+:12]), .o_data(C[50][2]), .i_clk(i_clk));
Mul0000000001  u_0000000262_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[818*12+:12]), .o_data(A[50][3]), .i_clk(i_clk));
Mul0000000001  u_0000000263_Mul0000000001(.i_data_1(c_plus_d[50][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[50][3]), .i_clk(i_clk));
Mul0000000001  u_0000000264_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[818*12+:12]), .o_data(C[50][3]), .i_clk(i_clk));
Mul0000000001  u_0000000265_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[51*12+:12]), .o_data(A[51][0]), .i_clk(i_clk));
Mul0000000001  u_0000000266_Mul0000000001(.i_data_1(c_plus_d[51][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[51][0]), .i_clk(i_clk));
Mul0000000001  u_0000000267_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[51*12+:12]), .o_data(C[51][0]), .i_clk(i_clk));
Mul0000000001  u_0000000268_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[307*12+:12]), .o_data(A[51][1]), .i_clk(i_clk));
Mul0000000001  u_0000000269_Mul0000000001(.i_data_1(c_plus_d[51][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[51][1]), .i_clk(i_clk));
Mul0000000001  u_000000026A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[307*12+:12]), .o_data(C[51][1]), .i_clk(i_clk));
Mul0000000001  u_000000026B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[563*12+:12]), .o_data(A[51][2]), .i_clk(i_clk));
Mul0000000001  u_000000026C_Mul0000000001(.i_data_1(c_plus_d[51][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[51][2]), .i_clk(i_clk));
Mul0000000001  u_000000026D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[563*12+:12]), .o_data(C[51][2]), .i_clk(i_clk));
Mul0000000001  u_000000026E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[819*12+:12]), .o_data(A[51][3]), .i_clk(i_clk));
Mul0000000001  u_000000026F_Mul0000000001(.i_data_1(c_plus_d[51][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[51][3]), .i_clk(i_clk));
Mul0000000001  u_0000000270_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[819*12+:12]), .o_data(C[51][3]), .i_clk(i_clk));
Mul0000000001  u_0000000271_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[52*12+:12]), .o_data(A[52][0]), .i_clk(i_clk));
Mul0000000001  u_0000000272_Mul0000000001(.i_data_1(c_plus_d[52][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[52][0]), .i_clk(i_clk));
Mul0000000001  u_0000000273_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[52*12+:12]), .o_data(C[52][0]), .i_clk(i_clk));
Mul0000000001  u_0000000274_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[308*12+:12]), .o_data(A[52][1]), .i_clk(i_clk));
Mul0000000001  u_0000000275_Mul0000000001(.i_data_1(c_plus_d[52][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[52][1]), .i_clk(i_clk));
Mul0000000001  u_0000000276_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[308*12+:12]), .o_data(C[52][1]), .i_clk(i_clk));
Mul0000000001  u_0000000277_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[564*12+:12]), .o_data(A[52][2]), .i_clk(i_clk));
Mul0000000001  u_0000000278_Mul0000000001(.i_data_1(c_plus_d[52][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[52][2]), .i_clk(i_clk));
Mul0000000001  u_0000000279_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[564*12+:12]), .o_data(C[52][2]), .i_clk(i_clk));
Mul0000000001  u_000000027A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[820*12+:12]), .o_data(A[52][3]), .i_clk(i_clk));
Mul0000000001  u_000000027B_Mul0000000001(.i_data_1(c_plus_d[52][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[52][3]), .i_clk(i_clk));
Mul0000000001  u_000000027C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[820*12+:12]), .o_data(C[52][3]), .i_clk(i_clk));
Mul0000000001  u_000000027D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[53*12+:12]), .o_data(A[53][0]), .i_clk(i_clk));
Mul0000000001  u_000000027E_Mul0000000001(.i_data_1(c_plus_d[53][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[53][0]), .i_clk(i_clk));
Mul0000000001  u_000000027F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[53*12+:12]), .o_data(C[53][0]), .i_clk(i_clk));
Mul0000000001  u_0000000280_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[309*12+:12]), .o_data(A[53][1]), .i_clk(i_clk));
Mul0000000001  u_0000000281_Mul0000000001(.i_data_1(c_plus_d[53][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[53][1]), .i_clk(i_clk));
Mul0000000001  u_0000000282_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[309*12+:12]), .o_data(C[53][1]), .i_clk(i_clk));
Mul0000000001  u_0000000283_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[565*12+:12]), .o_data(A[53][2]), .i_clk(i_clk));
Mul0000000001  u_0000000284_Mul0000000001(.i_data_1(c_plus_d[53][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[53][2]), .i_clk(i_clk));
Mul0000000001  u_0000000285_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[565*12+:12]), .o_data(C[53][2]), .i_clk(i_clk));
Mul0000000001  u_0000000286_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[821*12+:12]), .o_data(A[53][3]), .i_clk(i_clk));
Mul0000000001  u_0000000287_Mul0000000001(.i_data_1(c_plus_d[53][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[53][3]), .i_clk(i_clk));
Mul0000000001  u_0000000288_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[821*12+:12]), .o_data(C[53][3]), .i_clk(i_clk));
Mul0000000001  u_0000000289_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[54*12+:12]), .o_data(A[54][0]), .i_clk(i_clk));
Mul0000000001  u_000000028A_Mul0000000001(.i_data_1(c_plus_d[54][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[54][0]), .i_clk(i_clk));
Mul0000000001  u_000000028B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[54*12+:12]), .o_data(C[54][0]), .i_clk(i_clk));
Mul0000000001  u_000000028C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[310*12+:12]), .o_data(A[54][1]), .i_clk(i_clk));
Mul0000000001  u_000000028D_Mul0000000001(.i_data_1(c_plus_d[54][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[54][1]), .i_clk(i_clk));
Mul0000000001  u_000000028E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[310*12+:12]), .o_data(C[54][1]), .i_clk(i_clk));
Mul0000000001  u_000000028F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[566*12+:12]), .o_data(A[54][2]), .i_clk(i_clk));
Mul0000000001  u_0000000290_Mul0000000001(.i_data_1(c_plus_d[54][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[54][2]), .i_clk(i_clk));
Mul0000000001  u_0000000291_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[566*12+:12]), .o_data(C[54][2]), .i_clk(i_clk));
Mul0000000001  u_0000000292_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[822*12+:12]), .o_data(A[54][3]), .i_clk(i_clk));
Mul0000000001  u_0000000293_Mul0000000001(.i_data_1(c_plus_d[54][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[54][3]), .i_clk(i_clk));
Mul0000000001  u_0000000294_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[822*12+:12]), .o_data(C[54][3]), .i_clk(i_clk));
Mul0000000001  u_0000000295_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[55*12+:12]), .o_data(A[55][0]), .i_clk(i_clk));
Mul0000000001  u_0000000296_Mul0000000001(.i_data_1(c_plus_d[55][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[55][0]), .i_clk(i_clk));
Mul0000000001  u_0000000297_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[55*12+:12]), .o_data(C[55][0]), .i_clk(i_clk));
Mul0000000001  u_0000000298_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[311*12+:12]), .o_data(A[55][1]), .i_clk(i_clk));
Mul0000000001  u_0000000299_Mul0000000001(.i_data_1(c_plus_d[55][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[55][1]), .i_clk(i_clk));
Mul0000000001  u_000000029A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[311*12+:12]), .o_data(C[55][1]), .i_clk(i_clk));
Mul0000000001  u_000000029B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[567*12+:12]), .o_data(A[55][2]), .i_clk(i_clk));
Mul0000000001  u_000000029C_Mul0000000001(.i_data_1(c_plus_d[55][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[55][2]), .i_clk(i_clk));
Mul0000000001  u_000000029D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[567*12+:12]), .o_data(C[55][2]), .i_clk(i_clk));
Mul0000000001  u_000000029E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[823*12+:12]), .o_data(A[55][3]), .i_clk(i_clk));
Mul0000000001  u_000000029F_Mul0000000001(.i_data_1(c_plus_d[55][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[55][3]), .i_clk(i_clk));
Mul0000000001  u_00000002A0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[823*12+:12]), .o_data(C[55][3]), .i_clk(i_clk));
Mul0000000001  u_00000002A1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[56*12+:12]), .o_data(A[56][0]), .i_clk(i_clk));
Mul0000000001  u_00000002A2_Mul0000000001(.i_data_1(c_plus_d[56][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[56][0]), .i_clk(i_clk));
Mul0000000001  u_00000002A3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[56*12+:12]), .o_data(C[56][0]), .i_clk(i_clk));
Mul0000000001  u_00000002A4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[312*12+:12]), .o_data(A[56][1]), .i_clk(i_clk));
Mul0000000001  u_00000002A5_Mul0000000001(.i_data_1(c_plus_d[56][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[56][1]), .i_clk(i_clk));
Mul0000000001  u_00000002A6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[312*12+:12]), .o_data(C[56][1]), .i_clk(i_clk));
Mul0000000001  u_00000002A7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[568*12+:12]), .o_data(A[56][2]), .i_clk(i_clk));
Mul0000000001  u_00000002A8_Mul0000000001(.i_data_1(c_plus_d[56][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[56][2]), .i_clk(i_clk));
Mul0000000001  u_00000002A9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[568*12+:12]), .o_data(C[56][2]), .i_clk(i_clk));
Mul0000000001  u_00000002AA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[824*12+:12]), .o_data(A[56][3]), .i_clk(i_clk));
Mul0000000001  u_00000002AB_Mul0000000001(.i_data_1(c_plus_d[56][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[56][3]), .i_clk(i_clk));
Mul0000000001  u_00000002AC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[824*12+:12]), .o_data(C[56][3]), .i_clk(i_clk));
Mul0000000001  u_00000002AD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[57*12+:12]), .o_data(A[57][0]), .i_clk(i_clk));
Mul0000000001  u_00000002AE_Mul0000000001(.i_data_1(c_plus_d[57][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[57][0]), .i_clk(i_clk));
Mul0000000001  u_00000002AF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[57*12+:12]), .o_data(C[57][0]), .i_clk(i_clk));
Mul0000000001  u_00000002B0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[313*12+:12]), .o_data(A[57][1]), .i_clk(i_clk));
Mul0000000001  u_00000002B1_Mul0000000001(.i_data_1(c_plus_d[57][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[57][1]), .i_clk(i_clk));
Mul0000000001  u_00000002B2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[313*12+:12]), .o_data(C[57][1]), .i_clk(i_clk));
Mul0000000001  u_00000002B3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[569*12+:12]), .o_data(A[57][2]), .i_clk(i_clk));
Mul0000000001  u_00000002B4_Mul0000000001(.i_data_1(c_plus_d[57][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[57][2]), .i_clk(i_clk));
Mul0000000001  u_00000002B5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[569*12+:12]), .o_data(C[57][2]), .i_clk(i_clk));
Mul0000000001  u_00000002B6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[825*12+:12]), .o_data(A[57][3]), .i_clk(i_clk));
Mul0000000001  u_00000002B7_Mul0000000001(.i_data_1(c_plus_d[57][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[57][3]), .i_clk(i_clk));
Mul0000000001  u_00000002B8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[825*12+:12]), .o_data(C[57][3]), .i_clk(i_clk));
Mul0000000001  u_00000002B9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[58*12+:12]), .o_data(A[58][0]), .i_clk(i_clk));
Mul0000000001  u_00000002BA_Mul0000000001(.i_data_1(c_plus_d[58][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[58][0]), .i_clk(i_clk));
Mul0000000001  u_00000002BB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[58*12+:12]), .o_data(C[58][0]), .i_clk(i_clk));
Mul0000000001  u_00000002BC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[314*12+:12]), .o_data(A[58][1]), .i_clk(i_clk));
Mul0000000001  u_00000002BD_Mul0000000001(.i_data_1(c_plus_d[58][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[58][1]), .i_clk(i_clk));
Mul0000000001  u_00000002BE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[314*12+:12]), .o_data(C[58][1]), .i_clk(i_clk));
Mul0000000001  u_00000002BF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[570*12+:12]), .o_data(A[58][2]), .i_clk(i_clk));
Mul0000000001  u_00000002C0_Mul0000000001(.i_data_1(c_plus_d[58][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[58][2]), .i_clk(i_clk));
Mul0000000001  u_00000002C1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[570*12+:12]), .o_data(C[58][2]), .i_clk(i_clk));
Mul0000000001  u_00000002C2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[826*12+:12]), .o_data(A[58][3]), .i_clk(i_clk));
Mul0000000001  u_00000002C3_Mul0000000001(.i_data_1(c_plus_d[58][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[58][3]), .i_clk(i_clk));
Mul0000000001  u_00000002C4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[826*12+:12]), .o_data(C[58][3]), .i_clk(i_clk));
Mul0000000001  u_00000002C5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[59*12+:12]), .o_data(A[59][0]), .i_clk(i_clk));
Mul0000000001  u_00000002C6_Mul0000000001(.i_data_1(c_plus_d[59][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[59][0]), .i_clk(i_clk));
Mul0000000001  u_00000002C7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[59*12+:12]), .o_data(C[59][0]), .i_clk(i_clk));
Mul0000000001  u_00000002C8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[315*12+:12]), .o_data(A[59][1]), .i_clk(i_clk));
Mul0000000001  u_00000002C9_Mul0000000001(.i_data_1(c_plus_d[59][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[59][1]), .i_clk(i_clk));
Mul0000000001  u_00000002CA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[315*12+:12]), .o_data(C[59][1]), .i_clk(i_clk));
Mul0000000001  u_00000002CB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[571*12+:12]), .o_data(A[59][2]), .i_clk(i_clk));
Mul0000000001  u_00000002CC_Mul0000000001(.i_data_1(c_plus_d[59][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[59][2]), .i_clk(i_clk));
Mul0000000001  u_00000002CD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[571*12+:12]), .o_data(C[59][2]), .i_clk(i_clk));
Mul0000000001  u_00000002CE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[827*12+:12]), .o_data(A[59][3]), .i_clk(i_clk));
Mul0000000001  u_00000002CF_Mul0000000001(.i_data_1(c_plus_d[59][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[59][3]), .i_clk(i_clk));
Mul0000000001  u_00000002D0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[827*12+:12]), .o_data(C[59][3]), .i_clk(i_clk));
Mul0000000001  u_00000002D1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[60*12+:12]), .o_data(A[60][0]), .i_clk(i_clk));
Mul0000000001  u_00000002D2_Mul0000000001(.i_data_1(c_plus_d[60][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[60][0]), .i_clk(i_clk));
Mul0000000001  u_00000002D3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[60*12+:12]), .o_data(C[60][0]), .i_clk(i_clk));
Mul0000000001  u_00000002D4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[316*12+:12]), .o_data(A[60][1]), .i_clk(i_clk));
Mul0000000001  u_00000002D5_Mul0000000001(.i_data_1(c_plus_d[60][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[60][1]), .i_clk(i_clk));
Mul0000000001  u_00000002D6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[316*12+:12]), .o_data(C[60][1]), .i_clk(i_clk));
Mul0000000001  u_00000002D7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[572*12+:12]), .o_data(A[60][2]), .i_clk(i_clk));
Mul0000000001  u_00000002D8_Mul0000000001(.i_data_1(c_plus_d[60][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[60][2]), .i_clk(i_clk));
Mul0000000001  u_00000002D9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[572*12+:12]), .o_data(C[60][2]), .i_clk(i_clk));
Mul0000000001  u_00000002DA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[828*12+:12]), .o_data(A[60][3]), .i_clk(i_clk));
Mul0000000001  u_00000002DB_Mul0000000001(.i_data_1(c_plus_d[60][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[60][3]), .i_clk(i_clk));
Mul0000000001  u_00000002DC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[828*12+:12]), .o_data(C[60][3]), .i_clk(i_clk));
Mul0000000001  u_00000002DD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[61*12+:12]), .o_data(A[61][0]), .i_clk(i_clk));
Mul0000000001  u_00000002DE_Mul0000000001(.i_data_1(c_plus_d[61][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[61][0]), .i_clk(i_clk));
Mul0000000001  u_00000002DF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[61*12+:12]), .o_data(C[61][0]), .i_clk(i_clk));
Mul0000000001  u_00000002E0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[317*12+:12]), .o_data(A[61][1]), .i_clk(i_clk));
Mul0000000001  u_00000002E1_Mul0000000001(.i_data_1(c_plus_d[61][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[61][1]), .i_clk(i_clk));
Mul0000000001  u_00000002E2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[317*12+:12]), .o_data(C[61][1]), .i_clk(i_clk));
Mul0000000001  u_00000002E3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[573*12+:12]), .o_data(A[61][2]), .i_clk(i_clk));
Mul0000000001  u_00000002E4_Mul0000000001(.i_data_1(c_plus_d[61][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[61][2]), .i_clk(i_clk));
Mul0000000001  u_00000002E5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[573*12+:12]), .o_data(C[61][2]), .i_clk(i_clk));
Mul0000000001  u_00000002E6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[829*12+:12]), .o_data(A[61][3]), .i_clk(i_clk));
Mul0000000001  u_00000002E7_Mul0000000001(.i_data_1(c_plus_d[61][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[61][3]), .i_clk(i_clk));
Mul0000000001  u_00000002E8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[829*12+:12]), .o_data(C[61][3]), .i_clk(i_clk));
Mul0000000001  u_00000002E9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[62*12+:12]), .o_data(A[62][0]), .i_clk(i_clk));
Mul0000000001  u_00000002EA_Mul0000000001(.i_data_1(c_plus_d[62][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[62][0]), .i_clk(i_clk));
Mul0000000001  u_00000002EB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[62*12+:12]), .o_data(C[62][0]), .i_clk(i_clk));
Mul0000000001  u_00000002EC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[318*12+:12]), .o_data(A[62][1]), .i_clk(i_clk));
Mul0000000001  u_00000002ED_Mul0000000001(.i_data_1(c_plus_d[62][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[62][1]), .i_clk(i_clk));
Mul0000000001  u_00000002EE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[318*12+:12]), .o_data(C[62][1]), .i_clk(i_clk));
Mul0000000001  u_00000002EF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[574*12+:12]), .o_data(A[62][2]), .i_clk(i_clk));
Mul0000000001  u_00000002F0_Mul0000000001(.i_data_1(c_plus_d[62][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[62][2]), .i_clk(i_clk));
Mul0000000001  u_00000002F1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[574*12+:12]), .o_data(C[62][2]), .i_clk(i_clk));
Mul0000000001  u_00000002F2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[830*12+:12]), .o_data(A[62][3]), .i_clk(i_clk));
Mul0000000001  u_00000002F3_Mul0000000001(.i_data_1(c_plus_d[62][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[62][3]), .i_clk(i_clk));
Mul0000000001  u_00000002F4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[830*12+:12]), .o_data(C[62][3]), .i_clk(i_clk));
Mul0000000001  u_00000002F5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[63*12+:12]), .o_data(A[63][0]), .i_clk(i_clk));
Mul0000000001  u_00000002F6_Mul0000000001(.i_data_1(c_plus_d[63][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[63][0]), .i_clk(i_clk));
Mul0000000001  u_00000002F7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[63*12+:12]), .o_data(C[63][0]), .i_clk(i_clk));
Mul0000000001  u_00000002F8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[319*12+:12]), .o_data(A[63][1]), .i_clk(i_clk));
Mul0000000001  u_00000002F9_Mul0000000001(.i_data_1(c_plus_d[63][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[63][1]), .i_clk(i_clk));
Mul0000000001  u_00000002FA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[319*12+:12]), .o_data(C[63][1]), .i_clk(i_clk));
Mul0000000001  u_00000002FB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[575*12+:12]), .o_data(A[63][2]), .i_clk(i_clk));
Mul0000000001  u_00000002FC_Mul0000000001(.i_data_1(c_plus_d[63][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[63][2]), .i_clk(i_clk));
Mul0000000001  u_00000002FD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[575*12+:12]), .o_data(C[63][2]), .i_clk(i_clk));
Mul0000000001  u_00000002FE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[831*12+:12]), .o_data(A[63][3]), .i_clk(i_clk));
Mul0000000001  u_00000002FF_Mul0000000001(.i_data_1(c_plus_d[63][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[63][3]), .i_clk(i_clk));
Mul0000000001  u_0000000300_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[831*12+:12]), .o_data(C[63][3]), .i_clk(i_clk));
Mul0000000001  u_0000000301_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[64*12+:12]), .o_data(A[64][0]), .i_clk(i_clk));
Mul0000000001  u_0000000302_Mul0000000001(.i_data_1(c_plus_d[64][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[64][0]), .i_clk(i_clk));
Mul0000000001  u_0000000303_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[64*12+:12]), .o_data(C[64][0]), .i_clk(i_clk));
Mul0000000001  u_0000000304_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[320*12+:12]), .o_data(A[64][1]), .i_clk(i_clk));
Mul0000000001  u_0000000305_Mul0000000001(.i_data_1(c_plus_d[64][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[64][1]), .i_clk(i_clk));
Mul0000000001  u_0000000306_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[320*12+:12]), .o_data(C[64][1]), .i_clk(i_clk));
Mul0000000001  u_0000000307_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[576*12+:12]), .o_data(A[64][2]), .i_clk(i_clk));
Mul0000000001  u_0000000308_Mul0000000001(.i_data_1(c_plus_d[64][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[64][2]), .i_clk(i_clk));
Mul0000000001  u_0000000309_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[576*12+:12]), .o_data(C[64][2]), .i_clk(i_clk));
Mul0000000001  u_000000030A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[832*12+:12]), .o_data(A[64][3]), .i_clk(i_clk));
Mul0000000001  u_000000030B_Mul0000000001(.i_data_1(c_plus_d[64][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[64][3]), .i_clk(i_clk));
Mul0000000001  u_000000030C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[832*12+:12]), .o_data(C[64][3]), .i_clk(i_clk));
Mul0000000001  u_000000030D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[65*12+:12]), .o_data(A[65][0]), .i_clk(i_clk));
Mul0000000001  u_000000030E_Mul0000000001(.i_data_1(c_plus_d[65][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[65][0]), .i_clk(i_clk));
Mul0000000001  u_000000030F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[65*12+:12]), .o_data(C[65][0]), .i_clk(i_clk));
Mul0000000001  u_0000000310_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[321*12+:12]), .o_data(A[65][1]), .i_clk(i_clk));
Mul0000000001  u_0000000311_Mul0000000001(.i_data_1(c_plus_d[65][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[65][1]), .i_clk(i_clk));
Mul0000000001  u_0000000312_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[321*12+:12]), .o_data(C[65][1]), .i_clk(i_clk));
Mul0000000001  u_0000000313_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[577*12+:12]), .o_data(A[65][2]), .i_clk(i_clk));
Mul0000000001  u_0000000314_Mul0000000001(.i_data_1(c_plus_d[65][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[65][2]), .i_clk(i_clk));
Mul0000000001  u_0000000315_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[577*12+:12]), .o_data(C[65][2]), .i_clk(i_clk));
Mul0000000001  u_0000000316_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[833*12+:12]), .o_data(A[65][3]), .i_clk(i_clk));
Mul0000000001  u_0000000317_Mul0000000001(.i_data_1(c_plus_d[65][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[65][3]), .i_clk(i_clk));
Mul0000000001  u_0000000318_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[833*12+:12]), .o_data(C[65][3]), .i_clk(i_clk));
Mul0000000001  u_0000000319_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[66*12+:12]), .o_data(A[66][0]), .i_clk(i_clk));
Mul0000000001  u_000000031A_Mul0000000001(.i_data_1(c_plus_d[66][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[66][0]), .i_clk(i_clk));
Mul0000000001  u_000000031B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[66*12+:12]), .o_data(C[66][0]), .i_clk(i_clk));
Mul0000000001  u_000000031C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[322*12+:12]), .o_data(A[66][1]), .i_clk(i_clk));
Mul0000000001  u_000000031D_Mul0000000001(.i_data_1(c_plus_d[66][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[66][1]), .i_clk(i_clk));
Mul0000000001  u_000000031E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[322*12+:12]), .o_data(C[66][1]), .i_clk(i_clk));
Mul0000000001  u_000000031F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[578*12+:12]), .o_data(A[66][2]), .i_clk(i_clk));
Mul0000000001  u_0000000320_Mul0000000001(.i_data_1(c_plus_d[66][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[66][2]), .i_clk(i_clk));
Mul0000000001  u_0000000321_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[578*12+:12]), .o_data(C[66][2]), .i_clk(i_clk));
Mul0000000001  u_0000000322_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[834*12+:12]), .o_data(A[66][3]), .i_clk(i_clk));
Mul0000000001  u_0000000323_Mul0000000001(.i_data_1(c_plus_d[66][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[66][3]), .i_clk(i_clk));
Mul0000000001  u_0000000324_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[834*12+:12]), .o_data(C[66][3]), .i_clk(i_clk));
Mul0000000001  u_0000000325_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[67*12+:12]), .o_data(A[67][0]), .i_clk(i_clk));
Mul0000000001  u_0000000326_Mul0000000001(.i_data_1(c_plus_d[67][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[67][0]), .i_clk(i_clk));
Mul0000000001  u_0000000327_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[67*12+:12]), .o_data(C[67][0]), .i_clk(i_clk));
Mul0000000001  u_0000000328_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[323*12+:12]), .o_data(A[67][1]), .i_clk(i_clk));
Mul0000000001  u_0000000329_Mul0000000001(.i_data_1(c_plus_d[67][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[67][1]), .i_clk(i_clk));
Mul0000000001  u_000000032A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[323*12+:12]), .o_data(C[67][1]), .i_clk(i_clk));
Mul0000000001  u_000000032B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[579*12+:12]), .o_data(A[67][2]), .i_clk(i_clk));
Mul0000000001  u_000000032C_Mul0000000001(.i_data_1(c_plus_d[67][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[67][2]), .i_clk(i_clk));
Mul0000000001  u_000000032D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[579*12+:12]), .o_data(C[67][2]), .i_clk(i_clk));
Mul0000000001  u_000000032E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[835*12+:12]), .o_data(A[67][3]), .i_clk(i_clk));
Mul0000000001  u_000000032F_Mul0000000001(.i_data_1(c_plus_d[67][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[67][3]), .i_clk(i_clk));
Mul0000000001  u_0000000330_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[835*12+:12]), .o_data(C[67][3]), .i_clk(i_clk));
Mul0000000001  u_0000000331_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[68*12+:12]), .o_data(A[68][0]), .i_clk(i_clk));
Mul0000000001  u_0000000332_Mul0000000001(.i_data_1(c_plus_d[68][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[68][0]), .i_clk(i_clk));
Mul0000000001  u_0000000333_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[68*12+:12]), .o_data(C[68][0]), .i_clk(i_clk));
Mul0000000001  u_0000000334_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[324*12+:12]), .o_data(A[68][1]), .i_clk(i_clk));
Mul0000000001  u_0000000335_Mul0000000001(.i_data_1(c_plus_d[68][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[68][1]), .i_clk(i_clk));
Mul0000000001  u_0000000336_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[324*12+:12]), .o_data(C[68][1]), .i_clk(i_clk));
Mul0000000001  u_0000000337_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[580*12+:12]), .o_data(A[68][2]), .i_clk(i_clk));
Mul0000000001  u_0000000338_Mul0000000001(.i_data_1(c_plus_d[68][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[68][2]), .i_clk(i_clk));
Mul0000000001  u_0000000339_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[580*12+:12]), .o_data(C[68][2]), .i_clk(i_clk));
Mul0000000001  u_000000033A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[836*12+:12]), .o_data(A[68][3]), .i_clk(i_clk));
Mul0000000001  u_000000033B_Mul0000000001(.i_data_1(c_plus_d[68][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[68][3]), .i_clk(i_clk));
Mul0000000001  u_000000033C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[836*12+:12]), .o_data(C[68][3]), .i_clk(i_clk));
Mul0000000001  u_000000033D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[69*12+:12]), .o_data(A[69][0]), .i_clk(i_clk));
Mul0000000001  u_000000033E_Mul0000000001(.i_data_1(c_plus_d[69][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[69][0]), .i_clk(i_clk));
Mul0000000001  u_000000033F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[69*12+:12]), .o_data(C[69][0]), .i_clk(i_clk));
Mul0000000001  u_0000000340_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[325*12+:12]), .o_data(A[69][1]), .i_clk(i_clk));
Mul0000000001  u_0000000341_Mul0000000001(.i_data_1(c_plus_d[69][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[69][1]), .i_clk(i_clk));
Mul0000000001  u_0000000342_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[325*12+:12]), .o_data(C[69][1]), .i_clk(i_clk));
Mul0000000001  u_0000000343_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[581*12+:12]), .o_data(A[69][2]), .i_clk(i_clk));
Mul0000000001  u_0000000344_Mul0000000001(.i_data_1(c_plus_d[69][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[69][2]), .i_clk(i_clk));
Mul0000000001  u_0000000345_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[581*12+:12]), .o_data(C[69][2]), .i_clk(i_clk));
Mul0000000001  u_0000000346_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[837*12+:12]), .o_data(A[69][3]), .i_clk(i_clk));
Mul0000000001  u_0000000347_Mul0000000001(.i_data_1(c_plus_d[69][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[69][3]), .i_clk(i_clk));
Mul0000000001  u_0000000348_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[837*12+:12]), .o_data(C[69][3]), .i_clk(i_clk));
Mul0000000001  u_0000000349_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[70*12+:12]), .o_data(A[70][0]), .i_clk(i_clk));
Mul0000000001  u_000000034A_Mul0000000001(.i_data_1(c_plus_d[70][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[70][0]), .i_clk(i_clk));
Mul0000000001  u_000000034B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[70*12+:12]), .o_data(C[70][0]), .i_clk(i_clk));
Mul0000000001  u_000000034C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[326*12+:12]), .o_data(A[70][1]), .i_clk(i_clk));
Mul0000000001  u_000000034D_Mul0000000001(.i_data_1(c_plus_d[70][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[70][1]), .i_clk(i_clk));
Mul0000000001  u_000000034E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[326*12+:12]), .o_data(C[70][1]), .i_clk(i_clk));
Mul0000000001  u_000000034F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[582*12+:12]), .o_data(A[70][2]), .i_clk(i_clk));
Mul0000000001  u_0000000350_Mul0000000001(.i_data_1(c_plus_d[70][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[70][2]), .i_clk(i_clk));
Mul0000000001  u_0000000351_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[582*12+:12]), .o_data(C[70][2]), .i_clk(i_clk));
Mul0000000001  u_0000000352_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[838*12+:12]), .o_data(A[70][3]), .i_clk(i_clk));
Mul0000000001  u_0000000353_Mul0000000001(.i_data_1(c_plus_d[70][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[70][3]), .i_clk(i_clk));
Mul0000000001  u_0000000354_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[838*12+:12]), .o_data(C[70][3]), .i_clk(i_clk));
Mul0000000001  u_0000000355_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[71*12+:12]), .o_data(A[71][0]), .i_clk(i_clk));
Mul0000000001  u_0000000356_Mul0000000001(.i_data_1(c_plus_d[71][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[71][0]), .i_clk(i_clk));
Mul0000000001  u_0000000357_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[71*12+:12]), .o_data(C[71][0]), .i_clk(i_clk));
Mul0000000001  u_0000000358_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[327*12+:12]), .o_data(A[71][1]), .i_clk(i_clk));
Mul0000000001  u_0000000359_Mul0000000001(.i_data_1(c_plus_d[71][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[71][1]), .i_clk(i_clk));
Mul0000000001  u_000000035A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[327*12+:12]), .o_data(C[71][1]), .i_clk(i_clk));
Mul0000000001  u_000000035B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[583*12+:12]), .o_data(A[71][2]), .i_clk(i_clk));
Mul0000000001  u_000000035C_Mul0000000001(.i_data_1(c_plus_d[71][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[71][2]), .i_clk(i_clk));
Mul0000000001  u_000000035D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[583*12+:12]), .o_data(C[71][2]), .i_clk(i_clk));
Mul0000000001  u_000000035E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[839*12+:12]), .o_data(A[71][3]), .i_clk(i_clk));
Mul0000000001  u_000000035F_Mul0000000001(.i_data_1(c_plus_d[71][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[71][3]), .i_clk(i_clk));
Mul0000000001  u_0000000360_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[839*12+:12]), .o_data(C[71][3]), .i_clk(i_clk));
Mul0000000001  u_0000000361_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[72*12+:12]), .o_data(A[72][0]), .i_clk(i_clk));
Mul0000000001  u_0000000362_Mul0000000001(.i_data_1(c_plus_d[72][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[72][0]), .i_clk(i_clk));
Mul0000000001  u_0000000363_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[72*12+:12]), .o_data(C[72][0]), .i_clk(i_clk));
Mul0000000001  u_0000000364_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[328*12+:12]), .o_data(A[72][1]), .i_clk(i_clk));
Mul0000000001  u_0000000365_Mul0000000001(.i_data_1(c_plus_d[72][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[72][1]), .i_clk(i_clk));
Mul0000000001  u_0000000366_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[328*12+:12]), .o_data(C[72][1]), .i_clk(i_clk));
Mul0000000001  u_0000000367_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[584*12+:12]), .o_data(A[72][2]), .i_clk(i_clk));
Mul0000000001  u_0000000368_Mul0000000001(.i_data_1(c_plus_d[72][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[72][2]), .i_clk(i_clk));
Mul0000000001  u_0000000369_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[584*12+:12]), .o_data(C[72][2]), .i_clk(i_clk));
Mul0000000001  u_000000036A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[840*12+:12]), .o_data(A[72][3]), .i_clk(i_clk));
Mul0000000001  u_000000036B_Mul0000000001(.i_data_1(c_plus_d[72][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[72][3]), .i_clk(i_clk));
Mul0000000001  u_000000036C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[840*12+:12]), .o_data(C[72][3]), .i_clk(i_clk));
Mul0000000001  u_000000036D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[73*12+:12]), .o_data(A[73][0]), .i_clk(i_clk));
Mul0000000001  u_000000036E_Mul0000000001(.i_data_1(c_plus_d[73][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[73][0]), .i_clk(i_clk));
Mul0000000001  u_000000036F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[73*12+:12]), .o_data(C[73][0]), .i_clk(i_clk));
Mul0000000001  u_0000000370_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[329*12+:12]), .o_data(A[73][1]), .i_clk(i_clk));
Mul0000000001  u_0000000371_Mul0000000001(.i_data_1(c_plus_d[73][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[73][1]), .i_clk(i_clk));
Mul0000000001  u_0000000372_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[329*12+:12]), .o_data(C[73][1]), .i_clk(i_clk));
Mul0000000001  u_0000000373_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[585*12+:12]), .o_data(A[73][2]), .i_clk(i_clk));
Mul0000000001  u_0000000374_Mul0000000001(.i_data_1(c_plus_d[73][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[73][2]), .i_clk(i_clk));
Mul0000000001  u_0000000375_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[585*12+:12]), .o_data(C[73][2]), .i_clk(i_clk));
Mul0000000001  u_0000000376_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[841*12+:12]), .o_data(A[73][3]), .i_clk(i_clk));
Mul0000000001  u_0000000377_Mul0000000001(.i_data_1(c_plus_d[73][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[73][3]), .i_clk(i_clk));
Mul0000000001  u_0000000378_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[841*12+:12]), .o_data(C[73][3]), .i_clk(i_clk));
Mul0000000001  u_0000000379_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[74*12+:12]), .o_data(A[74][0]), .i_clk(i_clk));
Mul0000000001  u_000000037A_Mul0000000001(.i_data_1(c_plus_d[74][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[74][0]), .i_clk(i_clk));
Mul0000000001  u_000000037B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[74*12+:12]), .o_data(C[74][0]), .i_clk(i_clk));
Mul0000000001  u_000000037C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[330*12+:12]), .o_data(A[74][1]), .i_clk(i_clk));
Mul0000000001  u_000000037D_Mul0000000001(.i_data_1(c_plus_d[74][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[74][1]), .i_clk(i_clk));
Mul0000000001  u_000000037E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[330*12+:12]), .o_data(C[74][1]), .i_clk(i_clk));
Mul0000000001  u_000000037F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[586*12+:12]), .o_data(A[74][2]), .i_clk(i_clk));
Mul0000000001  u_0000000380_Mul0000000001(.i_data_1(c_plus_d[74][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[74][2]), .i_clk(i_clk));
Mul0000000001  u_0000000381_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[586*12+:12]), .o_data(C[74][2]), .i_clk(i_clk));
Mul0000000001  u_0000000382_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[842*12+:12]), .o_data(A[74][3]), .i_clk(i_clk));
Mul0000000001  u_0000000383_Mul0000000001(.i_data_1(c_plus_d[74][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[74][3]), .i_clk(i_clk));
Mul0000000001  u_0000000384_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[842*12+:12]), .o_data(C[74][3]), .i_clk(i_clk));
Mul0000000001  u_0000000385_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[75*12+:12]), .o_data(A[75][0]), .i_clk(i_clk));
Mul0000000001  u_0000000386_Mul0000000001(.i_data_1(c_plus_d[75][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[75][0]), .i_clk(i_clk));
Mul0000000001  u_0000000387_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[75*12+:12]), .o_data(C[75][0]), .i_clk(i_clk));
Mul0000000001  u_0000000388_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[331*12+:12]), .o_data(A[75][1]), .i_clk(i_clk));
Mul0000000001  u_0000000389_Mul0000000001(.i_data_1(c_plus_d[75][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[75][1]), .i_clk(i_clk));
Mul0000000001  u_000000038A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[331*12+:12]), .o_data(C[75][1]), .i_clk(i_clk));
Mul0000000001  u_000000038B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[587*12+:12]), .o_data(A[75][2]), .i_clk(i_clk));
Mul0000000001  u_000000038C_Mul0000000001(.i_data_1(c_plus_d[75][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[75][2]), .i_clk(i_clk));
Mul0000000001  u_000000038D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[587*12+:12]), .o_data(C[75][2]), .i_clk(i_clk));
Mul0000000001  u_000000038E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[843*12+:12]), .o_data(A[75][3]), .i_clk(i_clk));
Mul0000000001  u_000000038F_Mul0000000001(.i_data_1(c_plus_d[75][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[75][3]), .i_clk(i_clk));
Mul0000000001  u_0000000390_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[843*12+:12]), .o_data(C[75][3]), .i_clk(i_clk));
Mul0000000001  u_0000000391_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[76*12+:12]), .o_data(A[76][0]), .i_clk(i_clk));
Mul0000000001  u_0000000392_Mul0000000001(.i_data_1(c_plus_d[76][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[76][0]), .i_clk(i_clk));
Mul0000000001  u_0000000393_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[76*12+:12]), .o_data(C[76][0]), .i_clk(i_clk));
Mul0000000001  u_0000000394_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[332*12+:12]), .o_data(A[76][1]), .i_clk(i_clk));
Mul0000000001  u_0000000395_Mul0000000001(.i_data_1(c_plus_d[76][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[76][1]), .i_clk(i_clk));
Mul0000000001  u_0000000396_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[332*12+:12]), .o_data(C[76][1]), .i_clk(i_clk));
Mul0000000001  u_0000000397_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[588*12+:12]), .o_data(A[76][2]), .i_clk(i_clk));
Mul0000000001  u_0000000398_Mul0000000001(.i_data_1(c_plus_d[76][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[76][2]), .i_clk(i_clk));
Mul0000000001  u_0000000399_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[588*12+:12]), .o_data(C[76][2]), .i_clk(i_clk));
Mul0000000001  u_000000039A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[844*12+:12]), .o_data(A[76][3]), .i_clk(i_clk));
Mul0000000001  u_000000039B_Mul0000000001(.i_data_1(c_plus_d[76][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[76][3]), .i_clk(i_clk));
Mul0000000001  u_000000039C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[844*12+:12]), .o_data(C[76][3]), .i_clk(i_clk));
Mul0000000001  u_000000039D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[77*12+:12]), .o_data(A[77][0]), .i_clk(i_clk));
Mul0000000001  u_000000039E_Mul0000000001(.i_data_1(c_plus_d[77][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[77][0]), .i_clk(i_clk));
Mul0000000001  u_000000039F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[77*12+:12]), .o_data(C[77][0]), .i_clk(i_clk));
Mul0000000001  u_00000003A0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[333*12+:12]), .o_data(A[77][1]), .i_clk(i_clk));
Mul0000000001  u_00000003A1_Mul0000000001(.i_data_1(c_plus_d[77][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[77][1]), .i_clk(i_clk));
Mul0000000001  u_00000003A2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[333*12+:12]), .o_data(C[77][1]), .i_clk(i_clk));
Mul0000000001  u_00000003A3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[589*12+:12]), .o_data(A[77][2]), .i_clk(i_clk));
Mul0000000001  u_00000003A4_Mul0000000001(.i_data_1(c_plus_d[77][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[77][2]), .i_clk(i_clk));
Mul0000000001  u_00000003A5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[589*12+:12]), .o_data(C[77][2]), .i_clk(i_clk));
Mul0000000001  u_00000003A6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[845*12+:12]), .o_data(A[77][3]), .i_clk(i_clk));
Mul0000000001  u_00000003A7_Mul0000000001(.i_data_1(c_plus_d[77][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[77][3]), .i_clk(i_clk));
Mul0000000001  u_00000003A8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[845*12+:12]), .o_data(C[77][3]), .i_clk(i_clk));
Mul0000000001  u_00000003A9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[78*12+:12]), .o_data(A[78][0]), .i_clk(i_clk));
Mul0000000001  u_00000003AA_Mul0000000001(.i_data_1(c_plus_d[78][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[78][0]), .i_clk(i_clk));
Mul0000000001  u_00000003AB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[78*12+:12]), .o_data(C[78][0]), .i_clk(i_clk));
Mul0000000001  u_00000003AC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[334*12+:12]), .o_data(A[78][1]), .i_clk(i_clk));
Mul0000000001  u_00000003AD_Mul0000000001(.i_data_1(c_plus_d[78][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[78][1]), .i_clk(i_clk));
Mul0000000001  u_00000003AE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[334*12+:12]), .o_data(C[78][1]), .i_clk(i_clk));
Mul0000000001  u_00000003AF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[590*12+:12]), .o_data(A[78][2]), .i_clk(i_clk));
Mul0000000001  u_00000003B0_Mul0000000001(.i_data_1(c_plus_d[78][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[78][2]), .i_clk(i_clk));
Mul0000000001  u_00000003B1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[590*12+:12]), .o_data(C[78][2]), .i_clk(i_clk));
Mul0000000001  u_00000003B2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[846*12+:12]), .o_data(A[78][3]), .i_clk(i_clk));
Mul0000000001  u_00000003B3_Mul0000000001(.i_data_1(c_plus_d[78][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[78][3]), .i_clk(i_clk));
Mul0000000001  u_00000003B4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[846*12+:12]), .o_data(C[78][3]), .i_clk(i_clk));
Mul0000000001  u_00000003B5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[79*12+:12]), .o_data(A[79][0]), .i_clk(i_clk));
Mul0000000001  u_00000003B6_Mul0000000001(.i_data_1(c_plus_d[79][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[79][0]), .i_clk(i_clk));
Mul0000000001  u_00000003B7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[79*12+:12]), .o_data(C[79][0]), .i_clk(i_clk));
Mul0000000001  u_00000003B8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[335*12+:12]), .o_data(A[79][1]), .i_clk(i_clk));
Mul0000000001  u_00000003B9_Mul0000000001(.i_data_1(c_plus_d[79][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[79][1]), .i_clk(i_clk));
Mul0000000001  u_00000003BA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[335*12+:12]), .o_data(C[79][1]), .i_clk(i_clk));
Mul0000000001  u_00000003BB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[591*12+:12]), .o_data(A[79][2]), .i_clk(i_clk));
Mul0000000001  u_00000003BC_Mul0000000001(.i_data_1(c_plus_d[79][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[79][2]), .i_clk(i_clk));
Mul0000000001  u_00000003BD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[591*12+:12]), .o_data(C[79][2]), .i_clk(i_clk));
Mul0000000001  u_00000003BE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[847*12+:12]), .o_data(A[79][3]), .i_clk(i_clk));
Mul0000000001  u_00000003BF_Mul0000000001(.i_data_1(c_plus_d[79][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[79][3]), .i_clk(i_clk));
Mul0000000001  u_00000003C0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[847*12+:12]), .o_data(C[79][3]), .i_clk(i_clk));
Mul0000000001  u_00000003C1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[80*12+:12]), .o_data(A[80][0]), .i_clk(i_clk));
Mul0000000001  u_00000003C2_Mul0000000001(.i_data_1(c_plus_d[80][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[80][0]), .i_clk(i_clk));
Mul0000000001  u_00000003C3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[80*12+:12]), .o_data(C[80][0]), .i_clk(i_clk));
Mul0000000001  u_00000003C4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[336*12+:12]), .o_data(A[80][1]), .i_clk(i_clk));
Mul0000000001  u_00000003C5_Mul0000000001(.i_data_1(c_plus_d[80][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[80][1]), .i_clk(i_clk));
Mul0000000001  u_00000003C6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[336*12+:12]), .o_data(C[80][1]), .i_clk(i_clk));
Mul0000000001  u_00000003C7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[592*12+:12]), .o_data(A[80][2]), .i_clk(i_clk));
Mul0000000001  u_00000003C8_Mul0000000001(.i_data_1(c_plus_d[80][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[80][2]), .i_clk(i_clk));
Mul0000000001  u_00000003C9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[592*12+:12]), .o_data(C[80][2]), .i_clk(i_clk));
Mul0000000001  u_00000003CA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[848*12+:12]), .o_data(A[80][3]), .i_clk(i_clk));
Mul0000000001  u_00000003CB_Mul0000000001(.i_data_1(c_plus_d[80][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[80][3]), .i_clk(i_clk));
Mul0000000001  u_00000003CC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[848*12+:12]), .o_data(C[80][3]), .i_clk(i_clk));
Mul0000000001  u_00000003CD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[81*12+:12]), .o_data(A[81][0]), .i_clk(i_clk));
Mul0000000001  u_00000003CE_Mul0000000001(.i_data_1(c_plus_d[81][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[81][0]), .i_clk(i_clk));
Mul0000000001  u_00000003CF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[81*12+:12]), .o_data(C[81][0]), .i_clk(i_clk));
Mul0000000001  u_00000003D0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[337*12+:12]), .o_data(A[81][1]), .i_clk(i_clk));
Mul0000000001  u_00000003D1_Mul0000000001(.i_data_1(c_plus_d[81][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[81][1]), .i_clk(i_clk));
Mul0000000001  u_00000003D2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[337*12+:12]), .o_data(C[81][1]), .i_clk(i_clk));
Mul0000000001  u_00000003D3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[593*12+:12]), .o_data(A[81][2]), .i_clk(i_clk));
Mul0000000001  u_00000003D4_Mul0000000001(.i_data_1(c_plus_d[81][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[81][2]), .i_clk(i_clk));
Mul0000000001  u_00000003D5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[593*12+:12]), .o_data(C[81][2]), .i_clk(i_clk));
Mul0000000001  u_00000003D6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[849*12+:12]), .o_data(A[81][3]), .i_clk(i_clk));
Mul0000000001  u_00000003D7_Mul0000000001(.i_data_1(c_plus_d[81][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[81][3]), .i_clk(i_clk));
Mul0000000001  u_00000003D8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[849*12+:12]), .o_data(C[81][3]), .i_clk(i_clk));
Mul0000000001  u_00000003D9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[82*12+:12]), .o_data(A[82][0]), .i_clk(i_clk));
Mul0000000001  u_00000003DA_Mul0000000001(.i_data_1(c_plus_d[82][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[82][0]), .i_clk(i_clk));
Mul0000000001  u_00000003DB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[82*12+:12]), .o_data(C[82][0]), .i_clk(i_clk));
Mul0000000001  u_00000003DC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[338*12+:12]), .o_data(A[82][1]), .i_clk(i_clk));
Mul0000000001  u_00000003DD_Mul0000000001(.i_data_1(c_plus_d[82][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[82][1]), .i_clk(i_clk));
Mul0000000001  u_00000003DE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[338*12+:12]), .o_data(C[82][1]), .i_clk(i_clk));
Mul0000000001  u_00000003DF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[594*12+:12]), .o_data(A[82][2]), .i_clk(i_clk));
Mul0000000001  u_00000003E0_Mul0000000001(.i_data_1(c_plus_d[82][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[82][2]), .i_clk(i_clk));
Mul0000000001  u_00000003E1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[594*12+:12]), .o_data(C[82][2]), .i_clk(i_clk));
Mul0000000001  u_00000003E2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[850*12+:12]), .o_data(A[82][3]), .i_clk(i_clk));
Mul0000000001  u_00000003E3_Mul0000000001(.i_data_1(c_plus_d[82][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[82][3]), .i_clk(i_clk));
Mul0000000001  u_00000003E4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[850*12+:12]), .o_data(C[82][3]), .i_clk(i_clk));
Mul0000000001  u_00000003E5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[83*12+:12]), .o_data(A[83][0]), .i_clk(i_clk));
Mul0000000001  u_00000003E6_Mul0000000001(.i_data_1(c_plus_d[83][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[83][0]), .i_clk(i_clk));
Mul0000000001  u_00000003E7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[83*12+:12]), .o_data(C[83][0]), .i_clk(i_clk));
Mul0000000001  u_00000003E8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[339*12+:12]), .o_data(A[83][1]), .i_clk(i_clk));
Mul0000000001  u_00000003E9_Mul0000000001(.i_data_1(c_plus_d[83][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[83][1]), .i_clk(i_clk));
Mul0000000001  u_00000003EA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[339*12+:12]), .o_data(C[83][1]), .i_clk(i_clk));
Mul0000000001  u_00000003EB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[595*12+:12]), .o_data(A[83][2]), .i_clk(i_clk));
Mul0000000001  u_00000003EC_Mul0000000001(.i_data_1(c_plus_d[83][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[83][2]), .i_clk(i_clk));
Mul0000000001  u_00000003ED_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[595*12+:12]), .o_data(C[83][2]), .i_clk(i_clk));
Mul0000000001  u_00000003EE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[851*12+:12]), .o_data(A[83][3]), .i_clk(i_clk));
Mul0000000001  u_00000003EF_Mul0000000001(.i_data_1(c_plus_d[83][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[83][3]), .i_clk(i_clk));
Mul0000000001  u_00000003F0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[851*12+:12]), .o_data(C[83][3]), .i_clk(i_clk));
Mul0000000001  u_00000003F1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[84*12+:12]), .o_data(A[84][0]), .i_clk(i_clk));
Mul0000000001  u_00000003F2_Mul0000000001(.i_data_1(c_plus_d[84][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[84][0]), .i_clk(i_clk));
Mul0000000001  u_00000003F3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[84*12+:12]), .o_data(C[84][0]), .i_clk(i_clk));
Mul0000000001  u_00000003F4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[340*12+:12]), .o_data(A[84][1]), .i_clk(i_clk));
Mul0000000001  u_00000003F5_Mul0000000001(.i_data_1(c_plus_d[84][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[84][1]), .i_clk(i_clk));
Mul0000000001  u_00000003F6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[340*12+:12]), .o_data(C[84][1]), .i_clk(i_clk));
Mul0000000001  u_00000003F7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[596*12+:12]), .o_data(A[84][2]), .i_clk(i_clk));
Mul0000000001  u_00000003F8_Mul0000000001(.i_data_1(c_plus_d[84][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[84][2]), .i_clk(i_clk));
Mul0000000001  u_00000003F9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[596*12+:12]), .o_data(C[84][2]), .i_clk(i_clk));
Mul0000000001  u_00000003FA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[852*12+:12]), .o_data(A[84][3]), .i_clk(i_clk));
Mul0000000001  u_00000003FB_Mul0000000001(.i_data_1(c_plus_d[84][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[84][3]), .i_clk(i_clk));
Mul0000000001  u_00000003FC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[852*12+:12]), .o_data(C[84][3]), .i_clk(i_clk));
Mul0000000001  u_00000003FD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[85*12+:12]), .o_data(A[85][0]), .i_clk(i_clk));
Mul0000000001  u_00000003FE_Mul0000000001(.i_data_1(c_plus_d[85][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[85][0]), .i_clk(i_clk));
Mul0000000001  u_00000003FF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[85*12+:12]), .o_data(C[85][0]), .i_clk(i_clk));
Mul0000000001  u_0000000400_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[341*12+:12]), .o_data(A[85][1]), .i_clk(i_clk));
Mul0000000001  u_0000000401_Mul0000000001(.i_data_1(c_plus_d[85][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[85][1]), .i_clk(i_clk));
Mul0000000001  u_0000000402_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[341*12+:12]), .o_data(C[85][1]), .i_clk(i_clk));
Mul0000000001  u_0000000403_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[597*12+:12]), .o_data(A[85][2]), .i_clk(i_clk));
Mul0000000001  u_0000000404_Mul0000000001(.i_data_1(c_plus_d[85][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[85][2]), .i_clk(i_clk));
Mul0000000001  u_0000000405_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[597*12+:12]), .o_data(C[85][2]), .i_clk(i_clk));
Mul0000000001  u_0000000406_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[853*12+:12]), .o_data(A[85][3]), .i_clk(i_clk));
Mul0000000001  u_0000000407_Mul0000000001(.i_data_1(c_plus_d[85][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[85][3]), .i_clk(i_clk));
Mul0000000001  u_0000000408_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[853*12+:12]), .o_data(C[85][3]), .i_clk(i_clk));
Mul0000000001  u_0000000409_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[86*12+:12]), .o_data(A[86][0]), .i_clk(i_clk));
Mul0000000001  u_000000040A_Mul0000000001(.i_data_1(c_plus_d[86][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[86][0]), .i_clk(i_clk));
Mul0000000001  u_000000040B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[86*12+:12]), .o_data(C[86][0]), .i_clk(i_clk));
Mul0000000001  u_000000040C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[342*12+:12]), .o_data(A[86][1]), .i_clk(i_clk));
Mul0000000001  u_000000040D_Mul0000000001(.i_data_1(c_plus_d[86][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[86][1]), .i_clk(i_clk));
Mul0000000001  u_000000040E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[342*12+:12]), .o_data(C[86][1]), .i_clk(i_clk));
Mul0000000001  u_000000040F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[598*12+:12]), .o_data(A[86][2]), .i_clk(i_clk));
Mul0000000001  u_0000000410_Mul0000000001(.i_data_1(c_plus_d[86][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[86][2]), .i_clk(i_clk));
Mul0000000001  u_0000000411_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[598*12+:12]), .o_data(C[86][2]), .i_clk(i_clk));
Mul0000000001  u_0000000412_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[854*12+:12]), .o_data(A[86][3]), .i_clk(i_clk));
Mul0000000001  u_0000000413_Mul0000000001(.i_data_1(c_plus_d[86][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[86][3]), .i_clk(i_clk));
Mul0000000001  u_0000000414_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[854*12+:12]), .o_data(C[86][3]), .i_clk(i_clk));
Mul0000000001  u_0000000415_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[87*12+:12]), .o_data(A[87][0]), .i_clk(i_clk));
Mul0000000001  u_0000000416_Mul0000000001(.i_data_1(c_plus_d[87][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[87][0]), .i_clk(i_clk));
Mul0000000001  u_0000000417_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[87*12+:12]), .o_data(C[87][0]), .i_clk(i_clk));
Mul0000000001  u_0000000418_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[343*12+:12]), .o_data(A[87][1]), .i_clk(i_clk));
Mul0000000001  u_0000000419_Mul0000000001(.i_data_1(c_plus_d[87][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[87][1]), .i_clk(i_clk));
Mul0000000001  u_000000041A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[343*12+:12]), .o_data(C[87][1]), .i_clk(i_clk));
Mul0000000001  u_000000041B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[599*12+:12]), .o_data(A[87][2]), .i_clk(i_clk));
Mul0000000001  u_000000041C_Mul0000000001(.i_data_1(c_plus_d[87][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[87][2]), .i_clk(i_clk));
Mul0000000001  u_000000041D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[599*12+:12]), .o_data(C[87][2]), .i_clk(i_clk));
Mul0000000001  u_000000041E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[855*12+:12]), .o_data(A[87][3]), .i_clk(i_clk));
Mul0000000001  u_000000041F_Mul0000000001(.i_data_1(c_plus_d[87][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[87][3]), .i_clk(i_clk));
Mul0000000001  u_0000000420_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[855*12+:12]), .o_data(C[87][3]), .i_clk(i_clk));
Mul0000000001  u_0000000421_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[88*12+:12]), .o_data(A[88][0]), .i_clk(i_clk));
Mul0000000001  u_0000000422_Mul0000000001(.i_data_1(c_plus_d[88][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[88][0]), .i_clk(i_clk));
Mul0000000001  u_0000000423_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[88*12+:12]), .o_data(C[88][0]), .i_clk(i_clk));
Mul0000000001  u_0000000424_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[344*12+:12]), .o_data(A[88][1]), .i_clk(i_clk));
Mul0000000001  u_0000000425_Mul0000000001(.i_data_1(c_plus_d[88][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[88][1]), .i_clk(i_clk));
Mul0000000001  u_0000000426_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[344*12+:12]), .o_data(C[88][1]), .i_clk(i_clk));
Mul0000000001  u_0000000427_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[600*12+:12]), .o_data(A[88][2]), .i_clk(i_clk));
Mul0000000001  u_0000000428_Mul0000000001(.i_data_1(c_plus_d[88][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[88][2]), .i_clk(i_clk));
Mul0000000001  u_0000000429_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[600*12+:12]), .o_data(C[88][2]), .i_clk(i_clk));
Mul0000000001  u_000000042A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[856*12+:12]), .o_data(A[88][3]), .i_clk(i_clk));
Mul0000000001  u_000000042B_Mul0000000001(.i_data_1(c_plus_d[88][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[88][3]), .i_clk(i_clk));
Mul0000000001  u_000000042C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[856*12+:12]), .o_data(C[88][3]), .i_clk(i_clk));
Mul0000000001  u_000000042D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[89*12+:12]), .o_data(A[89][0]), .i_clk(i_clk));
Mul0000000001  u_000000042E_Mul0000000001(.i_data_1(c_plus_d[89][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[89][0]), .i_clk(i_clk));
Mul0000000001  u_000000042F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[89*12+:12]), .o_data(C[89][0]), .i_clk(i_clk));
Mul0000000001  u_0000000430_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[345*12+:12]), .o_data(A[89][1]), .i_clk(i_clk));
Mul0000000001  u_0000000431_Mul0000000001(.i_data_1(c_plus_d[89][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[89][1]), .i_clk(i_clk));
Mul0000000001  u_0000000432_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[345*12+:12]), .o_data(C[89][1]), .i_clk(i_clk));
Mul0000000001  u_0000000433_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[601*12+:12]), .o_data(A[89][2]), .i_clk(i_clk));
Mul0000000001  u_0000000434_Mul0000000001(.i_data_1(c_plus_d[89][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[89][2]), .i_clk(i_clk));
Mul0000000001  u_0000000435_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[601*12+:12]), .o_data(C[89][2]), .i_clk(i_clk));
Mul0000000001  u_0000000436_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[857*12+:12]), .o_data(A[89][3]), .i_clk(i_clk));
Mul0000000001  u_0000000437_Mul0000000001(.i_data_1(c_plus_d[89][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[89][3]), .i_clk(i_clk));
Mul0000000001  u_0000000438_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[857*12+:12]), .o_data(C[89][3]), .i_clk(i_clk));
Mul0000000001  u_0000000439_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[90*12+:12]), .o_data(A[90][0]), .i_clk(i_clk));
Mul0000000001  u_000000043A_Mul0000000001(.i_data_1(c_plus_d[90][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[90][0]), .i_clk(i_clk));
Mul0000000001  u_000000043B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[90*12+:12]), .o_data(C[90][0]), .i_clk(i_clk));
Mul0000000001  u_000000043C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[346*12+:12]), .o_data(A[90][1]), .i_clk(i_clk));
Mul0000000001  u_000000043D_Mul0000000001(.i_data_1(c_plus_d[90][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[90][1]), .i_clk(i_clk));
Mul0000000001  u_000000043E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[346*12+:12]), .o_data(C[90][1]), .i_clk(i_clk));
Mul0000000001  u_000000043F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[602*12+:12]), .o_data(A[90][2]), .i_clk(i_clk));
Mul0000000001  u_0000000440_Mul0000000001(.i_data_1(c_plus_d[90][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[90][2]), .i_clk(i_clk));
Mul0000000001  u_0000000441_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[602*12+:12]), .o_data(C[90][2]), .i_clk(i_clk));
Mul0000000001  u_0000000442_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[858*12+:12]), .o_data(A[90][3]), .i_clk(i_clk));
Mul0000000001  u_0000000443_Mul0000000001(.i_data_1(c_plus_d[90][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[90][3]), .i_clk(i_clk));
Mul0000000001  u_0000000444_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[858*12+:12]), .o_data(C[90][3]), .i_clk(i_clk));
Mul0000000001  u_0000000445_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[91*12+:12]), .o_data(A[91][0]), .i_clk(i_clk));
Mul0000000001  u_0000000446_Mul0000000001(.i_data_1(c_plus_d[91][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[91][0]), .i_clk(i_clk));
Mul0000000001  u_0000000447_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[91*12+:12]), .o_data(C[91][0]), .i_clk(i_clk));
Mul0000000001  u_0000000448_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[347*12+:12]), .o_data(A[91][1]), .i_clk(i_clk));
Mul0000000001  u_0000000449_Mul0000000001(.i_data_1(c_plus_d[91][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[91][1]), .i_clk(i_clk));
Mul0000000001  u_000000044A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[347*12+:12]), .o_data(C[91][1]), .i_clk(i_clk));
Mul0000000001  u_000000044B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[603*12+:12]), .o_data(A[91][2]), .i_clk(i_clk));
Mul0000000001  u_000000044C_Mul0000000001(.i_data_1(c_plus_d[91][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[91][2]), .i_clk(i_clk));
Mul0000000001  u_000000044D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[603*12+:12]), .o_data(C[91][2]), .i_clk(i_clk));
Mul0000000001  u_000000044E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[859*12+:12]), .o_data(A[91][3]), .i_clk(i_clk));
Mul0000000001  u_000000044F_Mul0000000001(.i_data_1(c_plus_d[91][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[91][3]), .i_clk(i_clk));
Mul0000000001  u_0000000450_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[859*12+:12]), .o_data(C[91][3]), .i_clk(i_clk));
Mul0000000001  u_0000000451_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[92*12+:12]), .o_data(A[92][0]), .i_clk(i_clk));
Mul0000000001  u_0000000452_Mul0000000001(.i_data_1(c_plus_d[92][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[92][0]), .i_clk(i_clk));
Mul0000000001  u_0000000453_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[92*12+:12]), .o_data(C[92][0]), .i_clk(i_clk));
Mul0000000001  u_0000000454_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[348*12+:12]), .o_data(A[92][1]), .i_clk(i_clk));
Mul0000000001  u_0000000455_Mul0000000001(.i_data_1(c_plus_d[92][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[92][1]), .i_clk(i_clk));
Mul0000000001  u_0000000456_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[348*12+:12]), .o_data(C[92][1]), .i_clk(i_clk));
Mul0000000001  u_0000000457_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[604*12+:12]), .o_data(A[92][2]), .i_clk(i_clk));
Mul0000000001  u_0000000458_Mul0000000001(.i_data_1(c_plus_d[92][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[92][2]), .i_clk(i_clk));
Mul0000000001  u_0000000459_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[604*12+:12]), .o_data(C[92][2]), .i_clk(i_clk));
Mul0000000001  u_000000045A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[860*12+:12]), .o_data(A[92][3]), .i_clk(i_clk));
Mul0000000001  u_000000045B_Mul0000000001(.i_data_1(c_plus_d[92][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[92][3]), .i_clk(i_clk));
Mul0000000001  u_000000045C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[860*12+:12]), .o_data(C[92][3]), .i_clk(i_clk));
Mul0000000001  u_000000045D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[93*12+:12]), .o_data(A[93][0]), .i_clk(i_clk));
Mul0000000001  u_000000045E_Mul0000000001(.i_data_1(c_plus_d[93][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[93][0]), .i_clk(i_clk));
Mul0000000001  u_000000045F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[93*12+:12]), .o_data(C[93][0]), .i_clk(i_clk));
Mul0000000001  u_0000000460_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[349*12+:12]), .o_data(A[93][1]), .i_clk(i_clk));
Mul0000000001  u_0000000461_Mul0000000001(.i_data_1(c_plus_d[93][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[93][1]), .i_clk(i_clk));
Mul0000000001  u_0000000462_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[349*12+:12]), .o_data(C[93][1]), .i_clk(i_clk));
Mul0000000001  u_0000000463_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[605*12+:12]), .o_data(A[93][2]), .i_clk(i_clk));
Mul0000000001  u_0000000464_Mul0000000001(.i_data_1(c_plus_d[93][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[93][2]), .i_clk(i_clk));
Mul0000000001  u_0000000465_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[605*12+:12]), .o_data(C[93][2]), .i_clk(i_clk));
Mul0000000001  u_0000000466_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[861*12+:12]), .o_data(A[93][3]), .i_clk(i_clk));
Mul0000000001  u_0000000467_Mul0000000001(.i_data_1(c_plus_d[93][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[93][3]), .i_clk(i_clk));
Mul0000000001  u_0000000468_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[861*12+:12]), .o_data(C[93][3]), .i_clk(i_clk));
Mul0000000001  u_0000000469_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[94*12+:12]), .o_data(A[94][0]), .i_clk(i_clk));
Mul0000000001  u_000000046A_Mul0000000001(.i_data_1(c_plus_d[94][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[94][0]), .i_clk(i_clk));
Mul0000000001  u_000000046B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[94*12+:12]), .o_data(C[94][0]), .i_clk(i_clk));
Mul0000000001  u_000000046C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[350*12+:12]), .o_data(A[94][1]), .i_clk(i_clk));
Mul0000000001  u_000000046D_Mul0000000001(.i_data_1(c_plus_d[94][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[94][1]), .i_clk(i_clk));
Mul0000000001  u_000000046E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[350*12+:12]), .o_data(C[94][1]), .i_clk(i_clk));
Mul0000000001  u_000000046F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[606*12+:12]), .o_data(A[94][2]), .i_clk(i_clk));
Mul0000000001  u_0000000470_Mul0000000001(.i_data_1(c_plus_d[94][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[94][2]), .i_clk(i_clk));
Mul0000000001  u_0000000471_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[606*12+:12]), .o_data(C[94][2]), .i_clk(i_clk));
Mul0000000001  u_0000000472_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[862*12+:12]), .o_data(A[94][3]), .i_clk(i_clk));
Mul0000000001  u_0000000473_Mul0000000001(.i_data_1(c_plus_d[94][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[94][3]), .i_clk(i_clk));
Mul0000000001  u_0000000474_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[862*12+:12]), .o_data(C[94][3]), .i_clk(i_clk));
Mul0000000001  u_0000000475_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[95*12+:12]), .o_data(A[95][0]), .i_clk(i_clk));
Mul0000000001  u_0000000476_Mul0000000001(.i_data_1(c_plus_d[95][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[95][0]), .i_clk(i_clk));
Mul0000000001  u_0000000477_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[95*12+:12]), .o_data(C[95][0]), .i_clk(i_clk));
Mul0000000001  u_0000000478_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[351*12+:12]), .o_data(A[95][1]), .i_clk(i_clk));
Mul0000000001  u_0000000479_Mul0000000001(.i_data_1(c_plus_d[95][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[95][1]), .i_clk(i_clk));
Mul0000000001  u_000000047A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[351*12+:12]), .o_data(C[95][1]), .i_clk(i_clk));
Mul0000000001  u_000000047B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[607*12+:12]), .o_data(A[95][2]), .i_clk(i_clk));
Mul0000000001  u_000000047C_Mul0000000001(.i_data_1(c_plus_d[95][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[95][2]), .i_clk(i_clk));
Mul0000000001  u_000000047D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[607*12+:12]), .o_data(C[95][2]), .i_clk(i_clk));
Mul0000000001  u_000000047E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[863*12+:12]), .o_data(A[95][3]), .i_clk(i_clk));
Mul0000000001  u_000000047F_Mul0000000001(.i_data_1(c_plus_d[95][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[95][3]), .i_clk(i_clk));
Mul0000000001  u_0000000480_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[863*12+:12]), .o_data(C[95][3]), .i_clk(i_clk));
Mul0000000001  u_0000000481_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[96*12+:12]), .o_data(A[96][0]), .i_clk(i_clk));
Mul0000000001  u_0000000482_Mul0000000001(.i_data_1(c_plus_d[96][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[96][0]), .i_clk(i_clk));
Mul0000000001  u_0000000483_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[96*12+:12]), .o_data(C[96][0]), .i_clk(i_clk));
Mul0000000001  u_0000000484_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[352*12+:12]), .o_data(A[96][1]), .i_clk(i_clk));
Mul0000000001  u_0000000485_Mul0000000001(.i_data_1(c_plus_d[96][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[96][1]), .i_clk(i_clk));
Mul0000000001  u_0000000486_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[352*12+:12]), .o_data(C[96][1]), .i_clk(i_clk));
Mul0000000001  u_0000000487_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[608*12+:12]), .o_data(A[96][2]), .i_clk(i_clk));
Mul0000000001  u_0000000488_Mul0000000001(.i_data_1(c_plus_d[96][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[96][2]), .i_clk(i_clk));
Mul0000000001  u_0000000489_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[608*12+:12]), .o_data(C[96][2]), .i_clk(i_clk));
Mul0000000001  u_000000048A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[864*12+:12]), .o_data(A[96][3]), .i_clk(i_clk));
Mul0000000001  u_000000048B_Mul0000000001(.i_data_1(c_plus_d[96][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[96][3]), .i_clk(i_clk));
Mul0000000001  u_000000048C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[864*12+:12]), .o_data(C[96][3]), .i_clk(i_clk));
Mul0000000001  u_000000048D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[97*12+:12]), .o_data(A[97][0]), .i_clk(i_clk));
Mul0000000001  u_000000048E_Mul0000000001(.i_data_1(c_plus_d[97][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[97][0]), .i_clk(i_clk));
Mul0000000001  u_000000048F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[97*12+:12]), .o_data(C[97][0]), .i_clk(i_clk));
Mul0000000001  u_0000000490_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[353*12+:12]), .o_data(A[97][1]), .i_clk(i_clk));
Mul0000000001  u_0000000491_Mul0000000001(.i_data_1(c_plus_d[97][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[97][1]), .i_clk(i_clk));
Mul0000000001  u_0000000492_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[353*12+:12]), .o_data(C[97][1]), .i_clk(i_clk));
Mul0000000001  u_0000000493_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[609*12+:12]), .o_data(A[97][2]), .i_clk(i_clk));
Mul0000000001  u_0000000494_Mul0000000001(.i_data_1(c_plus_d[97][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[97][2]), .i_clk(i_clk));
Mul0000000001  u_0000000495_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[609*12+:12]), .o_data(C[97][2]), .i_clk(i_clk));
Mul0000000001  u_0000000496_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[865*12+:12]), .o_data(A[97][3]), .i_clk(i_clk));
Mul0000000001  u_0000000497_Mul0000000001(.i_data_1(c_plus_d[97][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[97][3]), .i_clk(i_clk));
Mul0000000001  u_0000000498_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[865*12+:12]), .o_data(C[97][3]), .i_clk(i_clk));
Mul0000000001  u_0000000499_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[98*12+:12]), .o_data(A[98][0]), .i_clk(i_clk));
Mul0000000001  u_000000049A_Mul0000000001(.i_data_1(c_plus_d[98][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[98][0]), .i_clk(i_clk));
Mul0000000001  u_000000049B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[98*12+:12]), .o_data(C[98][0]), .i_clk(i_clk));
Mul0000000001  u_000000049C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[354*12+:12]), .o_data(A[98][1]), .i_clk(i_clk));
Mul0000000001  u_000000049D_Mul0000000001(.i_data_1(c_plus_d[98][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[98][1]), .i_clk(i_clk));
Mul0000000001  u_000000049E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[354*12+:12]), .o_data(C[98][1]), .i_clk(i_clk));
Mul0000000001  u_000000049F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[610*12+:12]), .o_data(A[98][2]), .i_clk(i_clk));
Mul0000000001  u_00000004A0_Mul0000000001(.i_data_1(c_plus_d[98][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[98][2]), .i_clk(i_clk));
Mul0000000001  u_00000004A1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[610*12+:12]), .o_data(C[98][2]), .i_clk(i_clk));
Mul0000000001  u_00000004A2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[866*12+:12]), .o_data(A[98][3]), .i_clk(i_clk));
Mul0000000001  u_00000004A3_Mul0000000001(.i_data_1(c_plus_d[98][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[98][3]), .i_clk(i_clk));
Mul0000000001  u_00000004A4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[866*12+:12]), .o_data(C[98][3]), .i_clk(i_clk));
Mul0000000001  u_00000004A5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[99*12+:12]), .o_data(A[99][0]), .i_clk(i_clk));
Mul0000000001  u_00000004A6_Mul0000000001(.i_data_1(c_plus_d[99][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[99][0]), .i_clk(i_clk));
Mul0000000001  u_00000004A7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[99*12+:12]), .o_data(C[99][0]), .i_clk(i_clk));
Mul0000000001  u_00000004A8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[355*12+:12]), .o_data(A[99][1]), .i_clk(i_clk));
Mul0000000001  u_00000004A9_Mul0000000001(.i_data_1(c_plus_d[99][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[99][1]), .i_clk(i_clk));
Mul0000000001  u_00000004AA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[355*12+:12]), .o_data(C[99][1]), .i_clk(i_clk));
Mul0000000001  u_00000004AB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[611*12+:12]), .o_data(A[99][2]), .i_clk(i_clk));
Mul0000000001  u_00000004AC_Mul0000000001(.i_data_1(c_plus_d[99][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[99][2]), .i_clk(i_clk));
Mul0000000001  u_00000004AD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[611*12+:12]), .o_data(C[99][2]), .i_clk(i_clk));
Mul0000000001  u_00000004AE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[867*12+:12]), .o_data(A[99][3]), .i_clk(i_clk));
Mul0000000001  u_00000004AF_Mul0000000001(.i_data_1(c_plus_d[99][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[99][3]), .i_clk(i_clk));
Mul0000000001  u_00000004B0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[867*12+:12]), .o_data(C[99][3]), .i_clk(i_clk));
Mul0000000001  u_00000004B1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[100*12+:12]), .o_data(A[100][0]), .i_clk(i_clk));
Mul0000000001  u_00000004B2_Mul0000000001(.i_data_1(c_plus_d[100][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[100][0]), .i_clk(i_clk));
Mul0000000001  u_00000004B3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[100*12+:12]), .o_data(C[100][0]), .i_clk(i_clk));
Mul0000000001  u_00000004B4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[356*12+:12]), .o_data(A[100][1]), .i_clk(i_clk));
Mul0000000001  u_00000004B5_Mul0000000001(.i_data_1(c_plus_d[100][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[100][1]), .i_clk(i_clk));
Mul0000000001  u_00000004B6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[356*12+:12]), .o_data(C[100][1]), .i_clk(i_clk));
Mul0000000001  u_00000004B7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[612*12+:12]), .o_data(A[100][2]), .i_clk(i_clk));
Mul0000000001  u_00000004B8_Mul0000000001(.i_data_1(c_plus_d[100][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[100][2]), .i_clk(i_clk));
Mul0000000001  u_00000004B9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[612*12+:12]), .o_data(C[100][2]), .i_clk(i_clk));
Mul0000000001  u_00000004BA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[868*12+:12]), .o_data(A[100][3]), .i_clk(i_clk));
Mul0000000001  u_00000004BB_Mul0000000001(.i_data_1(c_plus_d[100][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[100][3]), .i_clk(i_clk));
Mul0000000001  u_00000004BC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[868*12+:12]), .o_data(C[100][3]), .i_clk(i_clk));
Mul0000000001  u_00000004BD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[101*12+:12]), .o_data(A[101][0]), .i_clk(i_clk));
Mul0000000001  u_00000004BE_Mul0000000001(.i_data_1(c_plus_d[101][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[101][0]), .i_clk(i_clk));
Mul0000000001  u_00000004BF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[101*12+:12]), .o_data(C[101][0]), .i_clk(i_clk));
Mul0000000001  u_00000004C0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[357*12+:12]), .o_data(A[101][1]), .i_clk(i_clk));
Mul0000000001  u_00000004C1_Mul0000000001(.i_data_1(c_plus_d[101][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[101][1]), .i_clk(i_clk));
Mul0000000001  u_00000004C2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[357*12+:12]), .o_data(C[101][1]), .i_clk(i_clk));
Mul0000000001  u_00000004C3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[613*12+:12]), .o_data(A[101][2]), .i_clk(i_clk));
Mul0000000001  u_00000004C4_Mul0000000001(.i_data_1(c_plus_d[101][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[101][2]), .i_clk(i_clk));
Mul0000000001  u_00000004C5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[613*12+:12]), .o_data(C[101][2]), .i_clk(i_clk));
Mul0000000001  u_00000004C6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[869*12+:12]), .o_data(A[101][3]), .i_clk(i_clk));
Mul0000000001  u_00000004C7_Mul0000000001(.i_data_1(c_plus_d[101][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[101][3]), .i_clk(i_clk));
Mul0000000001  u_00000004C8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[869*12+:12]), .o_data(C[101][3]), .i_clk(i_clk));
Mul0000000001  u_00000004C9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[102*12+:12]), .o_data(A[102][0]), .i_clk(i_clk));
Mul0000000001  u_00000004CA_Mul0000000001(.i_data_1(c_plus_d[102][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[102][0]), .i_clk(i_clk));
Mul0000000001  u_00000004CB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[102*12+:12]), .o_data(C[102][0]), .i_clk(i_clk));
Mul0000000001  u_00000004CC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[358*12+:12]), .o_data(A[102][1]), .i_clk(i_clk));
Mul0000000001  u_00000004CD_Mul0000000001(.i_data_1(c_plus_d[102][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[102][1]), .i_clk(i_clk));
Mul0000000001  u_00000004CE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[358*12+:12]), .o_data(C[102][1]), .i_clk(i_clk));
Mul0000000001  u_00000004CF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[614*12+:12]), .o_data(A[102][2]), .i_clk(i_clk));
Mul0000000001  u_00000004D0_Mul0000000001(.i_data_1(c_plus_d[102][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[102][2]), .i_clk(i_clk));
Mul0000000001  u_00000004D1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[614*12+:12]), .o_data(C[102][2]), .i_clk(i_clk));
Mul0000000001  u_00000004D2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[870*12+:12]), .o_data(A[102][3]), .i_clk(i_clk));
Mul0000000001  u_00000004D3_Mul0000000001(.i_data_1(c_plus_d[102][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[102][3]), .i_clk(i_clk));
Mul0000000001  u_00000004D4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[870*12+:12]), .o_data(C[102][3]), .i_clk(i_clk));
Mul0000000001  u_00000004D5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[103*12+:12]), .o_data(A[103][0]), .i_clk(i_clk));
Mul0000000001  u_00000004D6_Mul0000000001(.i_data_1(c_plus_d[103][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[103][0]), .i_clk(i_clk));
Mul0000000001  u_00000004D7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[103*12+:12]), .o_data(C[103][0]), .i_clk(i_clk));
Mul0000000001  u_00000004D8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[359*12+:12]), .o_data(A[103][1]), .i_clk(i_clk));
Mul0000000001  u_00000004D9_Mul0000000001(.i_data_1(c_plus_d[103][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[103][1]), .i_clk(i_clk));
Mul0000000001  u_00000004DA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[359*12+:12]), .o_data(C[103][1]), .i_clk(i_clk));
Mul0000000001  u_00000004DB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[615*12+:12]), .o_data(A[103][2]), .i_clk(i_clk));
Mul0000000001  u_00000004DC_Mul0000000001(.i_data_1(c_plus_d[103][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[103][2]), .i_clk(i_clk));
Mul0000000001  u_00000004DD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[615*12+:12]), .o_data(C[103][2]), .i_clk(i_clk));
Mul0000000001  u_00000004DE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[871*12+:12]), .o_data(A[103][3]), .i_clk(i_clk));
Mul0000000001  u_00000004DF_Mul0000000001(.i_data_1(c_plus_d[103][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[103][3]), .i_clk(i_clk));
Mul0000000001  u_00000004E0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[871*12+:12]), .o_data(C[103][3]), .i_clk(i_clk));
Mul0000000001  u_00000004E1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[104*12+:12]), .o_data(A[104][0]), .i_clk(i_clk));
Mul0000000001  u_00000004E2_Mul0000000001(.i_data_1(c_plus_d[104][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[104][0]), .i_clk(i_clk));
Mul0000000001  u_00000004E3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[104*12+:12]), .o_data(C[104][0]), .i_clk(i_clk));
Mul0000000001  u_00000004E4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[360*12+:12]), .o_data(A[104][1]), .i_clk(i_clk));
Mul0000000001  u_00000004E5_Mul0000000001(.i_data_1(c_plus_d[104][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[104][1]), .i_clk(i_clk));
Mul0000000001  u_00000004E6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[360*12+:12]), .o_data(C[104][1]), .i_clk(i_clk));
Mul0000000001  u_00000004E7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[616*12+:12]), .o_data(A[104][2]), .i_clk(i_clk));
Mul0000000001  u_00000004E8_Mul0000000001(.i_data_1(c_plus_d[104][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[104][2]), .i_clk(i_clk));
Mul0000000001  u_00000004E9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[616*12+:12]), .o_data(C[104][2]), .i_clk(i_clk));
Mul0000000001  u_00000004EA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[872*12+:12]), .o_data(A[104][3]), .i_clk(i_clk));
Mul0000000001  u_00000004EB_Mul0000000001(.i_data_1(c_plus_d[104][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[104][3]), .i_clk(i_clk));
Mul0000000001  u_00000004EC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[872*12+:12]), .o_data(C[104][3]), .i_clk(i_clk));
Mul0000000001  u_00000004ED_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[105*12+:12]), .o_data(A[105][0]), .i_clk(i_clk));
Mul0000000001  u_00000004EE_Mul0000000001(.i_data_1(c_plus_d[105][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[105][0]), .i_clk(i_clk));
Mul0000000001  u_00000004EF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[105*12+:12]), .o_data(C[105][0]), .i_clk(i_clk));
Mul0000000001  u_00000004F0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[361*12+:12]), .o_data(A[105][1]), .i_clk(i_clk));
Mul0000000001  u_00000004F1_Mul0000000001(.i_data_1(c_plus_d[105][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[105][1]), .i_clk(i_clk));
Mul0000000001  u_00000004F2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[361*12+:12]), .o_data(C[105][1]), .i_clk(i_clk));
Mul0000000001  u_00000004F3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[617*12+:12]), .o_data(A[105][2]), .i_clk(i_clk));
Mul0000000001  u_00000004F4_Mul0000000001(.i_data_1(c_plus_d[105][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[105][2]), .i_clk(i_clk));
Mul0000000001  u_00000004F5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[617*12+:12]), .o_data(C[105][2]), .i_clk(i_clk));
Mul0000000001  u_00000004F6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[873*12+:12]), .o_data(A[105][3]), .i_clk(i_clk));
Mul0000000001  u_00000004F7_Mul0000000001(.i_data_1(c_plus_d[105][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[105][3]), .i_clk(i_clk));
Mul0000000001  u_00000004F8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[873*12+:12]), .o_data(C[105][3]), .i_clk(i_clk));
Mul0000000001  u_00000004F9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[106*12+:12]), .o_data(A[106][0]), .i_clk(i_clk));
Mul0000000001  u_00000004FA_Mul0000000001(.i_data_1(c_plus_d[106][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[106][0]), .i_clk(i_clk));
Mul0000000001  u_00000004FB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[106*12+:12]), .o_data(C[106][0]), .i_clk(i_clk));
Mul0000000001  u_00000004FC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[362*12+:12]), .o_data(A[106][1]), .i_clk(i_clk));
Mul0000000001  u_00000004FD_Mul0000000001(.i_data_1(c_plus_d[106][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[106][1]), .i_clk(i_clk));
Mul0000000001  u_00000004FE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[362*12+:12]), .o_data(C[106][1]), .i_clk(i_clk));
Mul0000000001  u_00000004FF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[618*12+:12]), .o_data(A[106][2]), .i_clk(i_clk));
Mul0000000001  u_0000000500_Mul0000000001(.i_data_1(c_plus_d[106][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[106][2]), .i_clk(i_clk));
Mul0000000001  u_0000000501_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[618*12+:12]), .o_data(C[106][2]), .i_clk(i_clk));
Mul0000000001  u_0000000502_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[874*12+:12]), .o_data(A[106][3]), .i_clk(i_clk));
Mul0000000001  u_0000000503_Mul0000000001(.i_data_1(c_plus_d[106][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[106][3]), .i_clk(i_clk));
Mul0000000001  u_0000000504_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[874*12+:12]), .o_data(C[106][3]), .i_clk(i_clk));
Mul0000000001  u_0000000505_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[107*12+:12]), .o_data(A[107][0]), .i_clk(i_clk));
Mul0000000001  u_0000000506_Mul0000000001(.i_data_1(c_plus_d[107][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[107][0]), .i_clk(i_clk));
Mul0000000001  u_0000000507_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[107*12+:12]), .o_data(C[107][0]), .i_clk(i_clk));
Mul0000000001  u_0000000508_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[363*12+:12]), .o_data(A[107][1]), .i_clk(i_clk));
Mul0000000001  u_0000000509_Mul0000000001(.i_data_1(c_plus_d[107][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[107][1]), .i_clk(i_clk));
Mul0000000001  u_000000050A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[363*12+:12]), .o_data(C[107][1]), .i_clk(i_clk));
Mul0000000001  u_000000050B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[619*12+:12]), .o_data(A[107][2]), .i_clk(i_clk));
Mul0000000001  u_000000050C_Mul0000000001(.i_data_1(c_plus_d[107][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[107][2]), .i_clk(i_clk));
Mul0000000001  u_000000050D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[619*12+:12]), .o_data(C[107][2]), .i_clk(i_clk));
Mul0000000001  u_000000050E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[875*12+:12]), .o_data(A[107][3]), .i_clk(i_clk));
Mul0000000001  u_000000050F_Mul0000000001(.i_data_1(c_plus_d[107][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[107][3]), .i_clk(i_clk));
Mul0000000001  u_0000000510_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[875*12+:12]), .o_data(C[107][3]), .i_clk(i_clk));
Mul0000000001  u_0000000511_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[108*12+:12]), .o_data(A[108][0]), .i_clk(i_clk));
Mul0000000001  u_0000000512_Mul0000000001(.i_data_1(c_plus_d[108][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[108][0]), .i_clk(i_clk));
Mul0000000001  u_0000000513_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[108*12+:12]), .o_data(C[108][0]), .i_clk(i_clk));
Mul0000000001  u_0000000514_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[364*12+:12]), .o_data(A[108][1]), .i_clk(i_clk));
Mul0000000001  u_0000000515_Mul0000000001(.i_data_1(c_plus_d[108][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[108][1]), .i_clk(i_clk));
Mul0000000001  u_0000000516_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[364*12+:12]), .o_data(C[108][1]), .i_clk(i_clk));
Mul0000000001  u_0000000517_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[620*12+:12]), .o_data(A[108][2]), .i_clk(i_clk));
Mul0000000001  u_0000000518_Mul0000000001(.i_data_1(c_plus_d[108][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[108][2]), .i_clk(i_clk));
Mul0000000001  u_0000000519_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[620*12+:12]), .o_data(C[108][2]), .i_clk(i_clk));
Mul0000000001  u_000000051A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[876*12+:12]), .o_data(A[108][3]), .i_clk(i_clk));
Mul0000000001  u_000000051B_Mul0000000001(.i_data_1(c_plus_d[108][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[108][3]), .i_clk(i_clk));
Mul0000000001  u_000000051C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[876*12+:12]), .o_data(C[108][3]), .i_clk(i_clk));
Mul0000000001  u_000000051D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[109*12+:12]), .o_data(A[109][0]), .i_clk(i_clk));
Mul0000000001  u_000000051E_Mul0000000001(.i_data_1(c_plus_d[109][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[109][0]), .i_clk(i_clk));
Mul0000000001  u_000000051F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[109*12+:12]), .o_data(C[109][0]), .i_clk(i_clk));
Mul0000000001  u_0000000520_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[365*12+:12]), .o_data(A[109][1]), .i_clk(i_clk));
Mul0000000001  u_0000000521_Mul0000000001(.i_data_1(c_plus_d[109][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[109][1]), .i_clk(i_clk));
Mul0000000001  u_0000000522_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[365*12+:12]), .o_data(C[109][1]), .i_clk(i_clk));
Mul0000000001  u_0000000523_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[621*12+:12]), .o_data(A[109][2]), .i_clk(i_clk));
Mul0000000001  u_0000000524_Mul0000000001(.i_data_1(c_plus_d[109][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[109][2]), .i_clk(i_clk));
Mul0000000001  u_0000000525_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[621*12+:12]), .o_data(C[109][2]), .i_clk(i_clk));
Mul0000000001  u_0000000526_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[877*12+:12]), .o_data(A[109][3]), .i_clk(i_clk));
Mul0000000001  u_0000000527_Mul0000000001(.i_data_1(c_plus_d[109][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[109][3]), .i_clk(i_clk));
Mul0000000001  u_0000000528_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[877*12+:12]), .o_data(C[109][3]), .i_clk(i_clk));
Mul0000000001  u_0000000529_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[110*12+:12]), .o_data(A[110][0]), .i_clk(i_clk));
Mul0000000001  u_000000052A_Mul0000000001(.i_data_1(c_plus_d[110][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[110][0]), .i_clk(i_clk));
Mul0000000001  u_000000052B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[110*12+:12]), .o_data(C[110][0]), .i_clk(i_clk));
Mul0000000001  u_000000052C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[366*12+:12]), .o_data(A[110][1]), .i_clk(i_clk));
Mul0000000001  u_000000052D_Mul0000000001(.i_data_1(c_plus_d[110][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[110][1]), .i_clk(i_clk));
Mul0000000001  u_000000052E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[366*12+:12]), .o_data(C[110][1]), .i_clk(i_clk));
Mul0000000001  u_000000052F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[622*12+:12]), .o_data(A[110][2]), .i_clk(i_clk));
Mul0000000001  u_0000000530_Mul0000000001(.i_data_1(c_plus_d[110][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[110][2]), .i_clk(i_clk));
Mul0000000001  u_0000000531_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[622*12+:12]), .o_data(C[110][2]), .i_clk(i_clk));
Mul0000000001  u_0000000532_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[878*12+:12]), .o_data(A[110][3]), .i_clk(i_clk));
Mul0000000001  u_0000000533_Mul0000000001(.i_data_1(c_plus_d[110][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[110][3]), .i_clk(i_clk));
Mul0000000001  u_0000000534_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[878*12+:12]), .o_data(C[110][3]), .i_clk(i_clk));
Mul0000000001  u_0000000535_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[111*12+:12]), .o_data(A[111][0]), .i_clk(i_clk));
Mul0000000001  u_0000000536_Mul0000000001(.i_data_1(c_plus_d[111][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[111][0]), .i_clk(i_clk));
Mul0000000001  u_0000000537_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[111*12+:12]), .o_data(C[111][0]), .i_clk(i_clk));
Mul0000000001  u_0000000538_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[367*12+:12]), .o_data(A[111][1]), .i_clk(i_clk));
Mul0000000001  u_0000000539_Mul0000000001(.i_data_1(c_plus_d[111][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[111][1]), .i_clk(i_clk));
Mul0000000001  u_000000053A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[367*12+:12]), .o_data(C[111][1]), .i_clk(i_clk));
Mul0000000001  u_000000053B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[623*12+:12]), .o_data(A[111][2]), .i_clk(i_clk));
Mul0000000001  u_000000053C_Mul0000000001(.i_data_1(c_plus_d[111][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[111][2]), .i_clk(i_clk));
Mul0000000001  u_000000053D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[623*12+:12]), .o_data(C[111][2]), .i_clk(i_clk));
Mul0000000001  u_000000053E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[879*12+:12]), .o_data(A[111][3]), .i_clk(i_clk));
Mul0000000001  u_000000053F_Mul0000000001(.i_data_1(c_plus_d[111][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[111][3]), .i_clk(i_clk));
Mul0000000001  u_0000000540_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[879*12+:12]), .o_data(C[111][3]), .i_clk(i_clk));
Mul0000000001  u_0000000541_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[112*12+:12]), .o_data(A[112][0]), .i_clk(i_clk));
Mul0000000001  u_0000000542_Mul0000000001(.i_data_1(c_plus_d[112][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[112][0]), .i_clk(i_clk));
Mul0000000001  u_0000000543_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[112*12+:12]), .o_data(C[112][0]), .i_clk(i_clk));
Mul0000000001  u_0000000544_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[368*12+:12]), .o_data(A[112][1]), .i_clk(i_clk));
Mul0000000001  u_0000000545_Mul0000000001(.i_data_1(c_plus_d[112][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[112][1]), .i_clk(i_clk));
Mul0000000001  u_0000000546_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[368*12+:12]), .o_data(C[112][1]), .i_clk(i_clk));
Mul0000000001  u_0000000547_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[624*12+:12]), .o_data(A[112][2]), .i_clk(i_clk));
Mul0000000001  u_0000000548_Mul0000000001(.i_data_1(c_plus_d[112][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[112][2]), .i_clk(i_clk));
Mul0000000001  u_0000000549_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[624*12+:12]), .o_data(C[112][2]), .i_clk(i_clk));
Mul0000000001  u_000000054A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[880*12+:12]), .o_data(A[112][3]), .i_clk(i_clk));
Mul0000000001  u_000000054B_Mul0000000001(.i_data_1(c_plus_d[112][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[112][3]), .i_clk(i_clk));
Mul0000000001  u_000000054C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[880*12+:12]), .o_data(C[112][3]), .i_clk(i_clk));
Mul0000000001  u_000000054D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[113*12+:12]), .o_data(A[113][0]), .i_clk(i_clk));
Mul0000000001  u_000000054E_Mul0000000001(.i_data_1(c_plus_d[113][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[113][0]), .i_clk(i_clk));
Mul0000000001  u_000000054F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[113*12+:12]), .o_data(C[113][0]), .i_clk(i_clk));
Mul0000000001  u_0000000550_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[369*12+:12]), .o_data(A[113][1]), .i_clk(i_clk));
Mul0000000001  u_0000000551_Mul0000000001(.i_data_1(c_plus_d[113][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[113][1]), .i_clk(i_clk));
Mul0000000001  u_0000000552_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[369*12+:12]), .o_data(C[113][1]), .i_clk(i_clk));
Mul0000000001  u_0000000553_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[625*12+:12]), .o_data(A[113][2]), .i_clk(i_clk));
Mul0000000001  u_0000000554_Mul0000000001(.i_data_1(c_plus_d[113][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[113][2]), .i_clk(i_clk));
Mul0000000001  u_0000000555_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[625*12+:12]), .o_data(C[113][2]), .i_clk(i_clk));
Mul0000000001  u_0000000556_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[881*12+:12]), .o_data(A[113][3]), .i_clk(i_clk));
Mul0000000001  u_0000000557_Mul0000000001(.i_data_1(c_plus_d[113][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[113][3]), .i_clk(i_clk));
Mul0000000001  u_0000000558_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[881*12+:12]), .o_data(C[113][3]), .i_clk(i_clk));
Mul0000000001  u_0000000559_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[114*12+:12]), .o_data(A[114][0]), .i_clk(i_clk));
Mul0000000001  u_000000055A_Mul0000000001(.i_data_1(c_plus_d[114][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[114][0]), .i_clk(i_clk));
Mul0000000001  u_000000055B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[114*12+:12]), .o_data(C[114][0]), .i_clk(i_clk));
Mul0000000001  u_000000055C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[370*12+:12]), .o_data(A[114][1]), .i_clk(i_clk));
Mul0000000001  u_000000055D_Mul0000000001(.i_data_1(c_plus_d[114][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[114][1]), .i_clk(i_clk));
Mul0000000001  u_000000055E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[370*12+:12]), .o_data(C[114][1]), .i_clk(i_clk));
Mul0000000001  u_000000055F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[626*12+:12]), .o_data(A[114][2]), .i_clk(i_clk));
Mul0000000001  u_0000000560_Mul0000000001(.i_data_1(c_plus_d[114][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[114][2]), .i_clk(i_clk));
Mul0000000001  u_0000000561_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[626*12+:12]), .o_data(C[114][2]), .i_clk(i_clk));
Mul0000000001  u_0000000562_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[882*12+:12]), .o_data(A[114][3]), .i_clk(i_clk));
Mul0000000001  u_0000000563_Mul0000000001(.i_data_1(c_plus_d[114][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[114][3]), .i_clk(i_clk));
Mul0000000001  u_0000000564_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[882*12+:12]), .o_data(C[114][3]), .i_clk(i_clk));
Mul0000000001  u_0000000565_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[115*12+:12]), .o_data(A[115][0]), .i_clk(i_clk));
Mul0000000001  u_0000000566_Mul0000000001(.i_data_1(c_plus_d[115][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[115][0]), .i_clk(i_clk));
Mul0000000001  u_0000000567_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[115*12+:12]), .o_data(C[115][0]), .i_clk(i_clk));
Mul0000000001  u_0000000568_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[371*12+:12]), .o_data(A[115][1]), .i_clk(i_clk));
Mul0000000001  u_0000000569_Mul0000000001(.i_data_1(c_plus_d[115][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[115][1]), .i_clk(i_clk));
Mul0000000001  u_000000056A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[371*12+:12]), .o_data(C[115][1]), .i_clk(i_clk));
Mul0000000001  u_000000056B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[627*12+:12]), .o_data(A[115][2]), .i_clk(i_clk));
Mul0000000001  u_000000056C_Mul0000000001(.i_data_1(c_plus_d[115][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[115][2]), .i_clk(i_clk));
Mul0000000001  u_000000056D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[627*12+:12]), .o_data(C[115][2]), .i_clk(i_clk));
Mul0000000001  u_000000056E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[883*12+:12]), .o_data(A[115][3]), .i_clk(i_clk));
Mul0000000001  u_000000056F_Mul0000000001(.i_data_1(c_plus_d[115][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[115][3]), .i_clk(i_clk));
Mul0000000001  u_0000000570_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[883*12+:12]), .o_data(C[115][3]), .i_clk(i_clk));
Mul0000000001  u_0000000571_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[116*12+:12]), .o_data(A[116][0]), .i_clk(i_clk));
Mul0000000001  u_0000000572_Mul0000000001(.i_data_1(c_plus_d[116][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[116][0]), .i_clk(i_clk));
Mul0000000001  u_0000000573_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[116*12+:12]), .o_data(C[116][0]), .i_clk(i_clk));
Mul0000000001  u_0000000574_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[372*12+:12]), .o_data(A[116][1]), .i_clk(i_clk));
Mul0000000001  u_0000000575_Mul0000000001(.i_data_1(c_plus_d[116][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[116][1]), .i_clk(i_clk));
Mul0000000001  u_0000000576_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[372*12+:12]), .o_data(C[116][1]), .i_clk(i_clk));
Mul0000000001  u_0000000577_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[628*12+:12]), .o_data(A[116][2]), .i_clk(i_clk));
Mul0000000001  u_0000000578_Mul0000000001(.i_data_1(c_plus_d[116][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[116][2]), .i_clk(i_clk));
Mul0000000001  u_0000000579_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[628*12+:12]), .o_data(C[116][2]), .i_clk(i_clk));
Mul0000000001  u_000000057A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[884*12+:12]), .o_data(A[116][3]), .i_clk(i_clk));
Mul0000000001  u_000000057B_Mul0000000001(.i_data_1(c_plus_d[116][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[116][3]), .i_clk(i_clk));
Mul0000000001  u_000000057C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[884*12+:12]), .o_data(C[116][3]), .i_clk(i_clk));
Mul0000000001  u_000000057D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[117*12+:12]), .o_data(A[117][0]), .i_clk(i_clk));
Mul0000000001  u_000000057E_Mul0000000001(.i_data_1(c_plus_d[117][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[117][0]), .i_clk(i_clk));
Mul0000000001  u_000000057F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[117*12+:12]), .o_data(C[117][0]), .i_clk(i_clk));
Mul0000000001  u_0000000580_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[373*12+:12]), .o_data(A[117][1]), .i_clk(i_clk));
Mul0000000001  u_0000000581_Mul0000000001(.i_data_1(c_plus_d[117][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[117][1]), .i_clk(i_clk));
Mul0000000001  u_0000000582_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[373*12+:12]), .o_data(C[117][1]), .i_clk(i_clk));
Mul0000000001  u_0000000583_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[629*12+:12]), .o_data(A[117][2]), .i_clk(i_clk));
Mul0000000001  u_0000000584_Mul0000000001(.i_data_1(c_plus_d[117][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[117][2]), .i_clk(i_clk));
Mul0000000001  u_0000000585_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[629*12+:12]), .o_data(C[117][2]), .i_clk(i_clk));
Mul0000000001  u_0000000586_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[885*12+:12]), .o_data(A[117][3]), .i_clk(i_clk));
Mul0000000001  u_0000000587_Mul0000000001(.i_data_1(c_plus_d[117][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[117][3]), .i_clk(i_clk));
Mul0000000001  u_0000000588_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[885*12+:12]), .o_data(C[117][3]), .i_clk(i_clk));
Mul0000000001  u_0000000589_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[118*12+:12]), .o_data(A[118][0]), .i_clk(i_clk));
Mul0000000001  u_000000058A_Mul0000000001(.i_data_1(c_plus_d[118][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[118][0]), .i_clk(i_clk));
Mul0000000001  u_000000058B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[118*12+:12]), .o_data(C[118][0]), .i_clk(i_clk));
Mul0000000001  u_000000058C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[374*12+:12]), .o_data(A[118][1]), .i_clk(i_clk));
Mul0000000001  u_000000058D_Mul0000000001(.i_data_1(c_plus_d[118][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[118][1]), .i_clk(i_clk));
Mul0000000001  u_000000058E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[374*12+:12]), .o_data(C[118][1]), .i_clk(i_clk));
Mul0000000001  u_000000058F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[630*12+:12]), .o_data(A[118][2]), .i_clk(i_clk));
Mul0000000001  u_0000000590_Mul0000000001(.i_data_1(c_plus_d[118][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[118][2]), .i_clk(i_clk));
Mul0000000001  u_0000000591_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[630*12+:12]), .o_data(C[118][2]), .i_clk(i_clk));
Mul0000000001  u_0000000592_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[886*12+:12]), .o_data(A[118][3]), .i_clk(i_clk));
Mul0000000001  u_0000000593_Mul0000000001(.i_data_1(c_plus_d[118][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[118][3]), .i_clk(i_clk));
Mul0000000001  u_0000000594_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[886*12+:12]), .o_data(C[118][3]), .i_clk(i_clk));
Mul0000000001  u_0000000595_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[119*12+:12]), .o_data(A[119][0]), .i_clk(i_clk));
Mul0000000001  u_0000000596_Mul0000000001(.i_data_1(c_plus_d[119][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[119][0]), .i_clk(i_clk));
Mul0000000001  u_0000000597_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[119*12+:12]), .o_data(C[119][0]), .i_clk(i_clk));
Mul0000000001  u_0000000598_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[375*12+:12]), .o_data(A[119][1]), .i_clk(i_clk));
Mul0000000001  u_0000000599_Mul0000000001(.i_data_1(c_plus_d[119][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[119][1]), .i_clk(i_clk));
Mul0000000001  u_000000059A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[375*12+:12]), .o_data(C[119][1]), .i_clk(i_clk));
Mul0000000001  u_000000059B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[631*12+:12]), .o_data(A[119][2]), .i_clk(i_clk));
Mul0000000001  u_000000059C_Mul0000000001(.i_data_1(c_plus_d[119][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[119][2]), .i_clk(i_clk));
Mul0000000001  u_000000059D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[631*12+:12]), .o_data(C[119][2]), .i_clk(i_clk));
Mul0000000001  u_000000059E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[887*12+:12]), .o_data(A[119][3]), .i_clk(i_clk));
Mul0000000001  u_000000059F_Mul0000000001(.i_data_1(c_plus_d[119][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[119][3]), .i_clk(i_clk));
Mul0000000001  u_00000005A0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[887*12+:12]), .o_data(C[119][3]), .i_clk(i_clk));
Mul0000000001  u_00000005A1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[120*12+:12]), .o_data(A[120][0]), .i_clk(i_clk));
Mul0000000001  u_00000005A2_Mul0000000001(.i_data_1(c_plus_d[120][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[120][0]), .i_clk(i_clk));
Mul0000000001  u_00000005A3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[120*12+:12]), .o_data(C[120][0]), .i_clk(i_clk));
Mul0000000001  u_00000005A4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[376*12+:12]), .o_data(A[120][1]), .i_clk(i_clk));
Mul0000000001  u_00000005A5_Mul0000000001(.i_data_1(c_plus_d[120][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[120][1]), .i_clk(i_clk));
Mul0000000001  u_00000005A6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[376*12+:12]), .o_data(C[120][1]), .i_clk(i_clk));
Mul0000000001  u_00000005A7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[632*12+:12]), .o_data(A[120][2]), .i_clk(i_clk));
Mul0000000001  u_00000005A8_Mul0000000001(.i_data_1(c_plus_d[120][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[120][2]), .i_clk(i_clk));
Mul0000000001  u_00000005A9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[632*12+:12]), .o_data(C[120][2]), .i_clk(i_clk));
Mul0000000001  u_00000005AA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[888*12+:12]), .o_data(A[120][3]), .i_clk(i_clk));
Mul0000000001  u_00000005AB_Mul0000000001(.i_data_1(c_plus_d[120][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[120][3]), .i_clk(i_clk));
Mul0000000001  u_00000005AC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[888*12+:12]), .o_data(C[120][3]), .i_clk(i_clk));
Mul0000000001  u_00000005AD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[121*12+:12]), .o_data(A[121][0]), .i_clk(i_clk));
Mul0000000001  u_00000005AE_Mul0000000001(.i_data_1(c_plus_d[121][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[121][0]), .i_clk(i_clk));
Mul0000000001  u_00000005AF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[121*12+:12]), .o_data(C[121][0]), .i_clk(i_clk));
Mul0000000001  u_00000005B0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[377*12+:12]), .o_data(A[121][1]), .i_clk(i_clk));
Mul0000000001  u_00000005B1_Mul0000000001(.i_data_1(c_plus_d[121][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[121][1]), .i_clk(i_clk));
Mul0000000001  u_00000005B2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[377*12+:12]), .o_data(C[121][1]), .i_clk(i_clk));
Mul0000000001  u_00000005B3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[633*12+:12]), .o_data(A[121][2]), .i_clk(i_clk));
Mul0000000001  u_00000005B4_Mul0000000001(.i_data_1(c_plus_d[121][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[121][2]), .i_clk(i_clk));
Mul0000000001  u_00000005B5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[633*12+:12]), .o_data(C[121][2]), .i_clk(i_clk));
Mul0000000001  u_00000005B6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[889*12+:12]), .o_data(A[121][3]), .i_clk(i_clk));
Mul0000000001  u_00000005B7_Mul0000000001(.i_data_1(c_plus_d[121][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[121][3]), .i_clk(i_clk));
Mul0000000001  u_00000005B8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[889*12+:12]), .o_data(C[121][3]), .i_clk(i_clk));
Mul0000000001  u_00000005B9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[122*12+:12]), .o_data(A[122][0]), .i_clk(i_clk));
Mul0000000001  u_00000005BA_Mul0000000001(.i_data_1(c_plus_d[122][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[122][0]), .i_clk(i_clk));
Mul0000000001  u_00000005BB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[122*12+:12]), .o_data(C[122][0]), .i_clk(i_clk));
Mul0000000001  u_00000005BC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[378*12+:12]), .o_data(A[122][1]), .i_clk(i_clk));
Mul0000000001  u_00000005BD_Mul0000000001(.i_data_1(c_plus_d[122][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[122][1]), .i_clk(i_clk));
Mul0000000001  u_00000005BE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[378*12+:12]), .o_data(C[122][1]), .i_clk(i_clk));
Mul0000000001  u_00000005BF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[634*12+:12]), .o_data(A[122][2]), .i_clk(i_clk));
Mul0000000001  u_00000005C0_Mul0000000001(.i_data_1(c_plus_d[122][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[122][2]), .i_clk(i_clk));
Mul0000000001  u_00000005C1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[634*12+:12]), .o_data(C[122][2]), .i_clk(i_clk));
Mul0000000001  u_00000005C2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[890*12+:12]), .o_data(A[122][3]), .i_clk(i_clk));
Mul0000000001  u_00000005C3_Mul0000000001(.i_data_1(c_plus_d[122][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[122][3]), .i_clk(i_clk));
Mul0000000001  u_00000005C4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[890*12+:12]), .o_data(C[122][3]), .i_clk(i_clk));
Mul0000000001  u_00000005C5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[123*12+:12]), .o_data(A[123][0]), .i_clk(i_clk));
Mul0000000001  u_00000005C6_Mul0000000001(.i_data_1(c_plus_d[123][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[123][0]), .i_clk(i_clk));
Mul0000000001  u_00000005C7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[123*12+:12]), .o_data(C[123][0]), .i_clk(i_clk));
Mul0000000001  u_00000005C8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[379*12+:12]), .o_data(A[123][1]), .i_clk(i_clk));
Mul0000000001  u_00000005C9_Mul0000000001(.i_data_1(c_plus_d[123][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[123][1]), .i_clk(i_clk));
Mul0000000001  u_00000005CA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[379*12+:12]), .o_data(C[123][1]), .i_clk(i_clk));
Mul0000000001  u_00000005CB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[635*12+:12]), .o_data(A[123][2]), .i_clk(i_clk));
Mul0000000001  u_00000005CC_Mul0000000001(.i_data_1(c_plus_d[123][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[123][2]), .i_clk(i_clk));
Mul0000000001  u_00000005CD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[635*12+:12]), .o_data(C[123][2]), .i_clk(i_clk));
Mul0000000001  u_00000005CE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[891*12+:12]), .o_data(A[123][3]), .i_clk(i_clk));
Mul0000000001  u_00000005CF_Mul0000000001(.i_data_1(c_plus_d[123][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[123][3]), .i_clk(i_clk));
Mul0000000001  u_00000005D0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[891*12+:12]), .o_data(C[123][3]), .i_clk(i_clk));
Mul0000000001  u_00000005D1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[124*12+:12]), .o_data(A[124][0]), .i_clk(i_clk));
Mul0000000001  u_00000005D2_Mul0000000001(.i_data_1(c_plus_d[124][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[124][0]), .i_clk(i_clk));
Mul0000000001  u_00000005D3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[124*12+:12]), .o_data(C[124][0]), .i_clk(i_clk));
Mul0000000001  u_00000005D4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[380*12+:12]), .o_data(A[124][1]), .i_clk(i_clk));
Mul0000000001  u_00000005D5_Mul0000000001(.i_data_1(c_plus_d[124][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[124][1]), .i_clk(i_clk));
Mul0000000001  u_00000005D6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[380*12+:12]), .o_data(C[124][1]), .i_clk(i_clk));
Mul0000000001  u_00000005D7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[636*12+:12]), .o_data(A[124][2]), .i_clk(i_clk));
Mul0000000001  u_00000005D8_Mul0000000001(.i_data_1(c_plus_d[124][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[124][2]), .i_clk(i_clk));
Mul0000000001  u_00000005D9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[636*12+:12]), .o_data(C[124][2]), .i_clk(i_clk));
Mul0000000001  u_00000005DA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[892*12+:12]), .o_data(A[124][3]), .i_clk(i_clk));
Mul0000000001  u_00000005DB_Mul0000000001(.i_data_1(c_plus_d[124][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[124][3]), .i_clk(i_clk));
Mul0000000001  u_00000005DC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[892*12+:12]), .o_data(C[124][3]), .i_clk(i_clk));
Mul0000000001  u_00000005DD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[125*12+:12]), .o_data(A[125][0]), .i_clk(i_clk));
Mul0000000001  u_00000005DE_Mul0000000001(.i_data_1(c_plus_d[125][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[125][0]), .i_clk(i_clk));
Mul0000000001  u_00000005DF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[125*12+:12]), .o_data(C[125][0]), .i_clk(i_clk));
Mul0000000001  u_00000005E0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[381*12+:12]), .o_data(A[125][1]), .i_clk(i_clk));
Mul0000000001  u_00000005E1_Mul0000000001(.i_data_1(c_plus_d[125][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[125][1]), .i_clk(i_clk));
Mul0000000001  u_00000005E2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[381*12+:12]), .o_data(C[125][1]), .i_clk(i_clk));
Mul0000000001  u_00000005E3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[637*12+:12]), .o_data(A[125][2]), .i_clk(i_clk));
Mul0000000001  u_00000005E4_Mul0000000001(.i_data_1(c_plus_d[125][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[125][2]), .i_clk(i_clk));
Mul0000000001  u_00000005E5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[637*12+:12]), .o_data(C[125][2]), .i_clk(i_clk));
Mul0000000001  u_00000005E6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[893*12+:12]), .o_data(A[125][3]), .i_clk(i_clk));
Mul0000000001  u_00000005E7_Mul0000000001(.i_data_1(c_plus_d[125][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[125][3]), .i_clk(i_clk));
Mul0000000001  u_00000005E8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[893*12+:12]), .o_data(C[125][3]), .i_clk(i_clk));
Mul0000000001  u_00000005E9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[126*12+:12]), .o_data(A[126][0]), .i_clk(i_clk));
Mul0000000001  u_00000005EA_Mul0000000001(.i_data_1(c_plus_d[126][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[126][0]), .i_clk(i_clk));
Mul0000000001  u_00000005EB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[126*12+:12]), .o_data(C[126][0]), .i_clk(i_clk));
Mul0000000001  u_00000005EC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[382*12+:12]), .o_data(A[126][1]), .i_clk(i_clk));
Mul0000000001  u_00000005ED_Mul0000000001(.i_data_1(c_plus_d[126][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[126][1]), .i_clk(i_clk));
Mul0000000001  u_00000005EE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[382*12+:12]), .o_data(C[126][1]), .i_clk(i_clk));
Mul0000000001  u_00000005EF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[638*12+:12]), .o_data(A[126][2]), .i_clk(i_clk));
Mul0000000001  u_00000005F0_Mul0000000001(.i_data_1(c_plus_d[126][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[126][2]), .i_clk(i_clk));
Mul0000000001  u_00000005F1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[638*12+:12]), .o_data(C[126][2]), .i_clk(i_clk));
Mul0000000001  u_00000005F2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[894*12+:12]), .o_data(A[126][3]), .i_clk(i_clk));
Mul0000000001  u_00000005F3_Mul0000000001(.i_data_1(c_plus_d[126][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[126][3]), .i_clk(i_clk));
Mul0000000001  u_00000005F4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[894*12+:12]), .o_data(C[126][3]), .i_clk(i_clk));
Mul0000000001  u_00000005F5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[127*12+:12]), .o_data(A[127][0]), .i_clk(i_clk));
Mul0000000001  u_00000005F6_Mul0000000001(.i_data_1(c_plus_d[127][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[127][0]), .i_clk(i_clk));
Mul0000000001  u_00000005F7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[127*12+:12]), .o_data(C[127][0]), .i_clk(i_clk));
Mul0000000001  u_00000005F8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[383*12+:12]), .o_data(A[127][1]), .i_clk(i_clk));
Mul0000000001  u_00000005F9_Mul0000000001(.i_data_1(c_plus_d[127][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[127][1]), .i_clk(i_clk));
Mul0000000001  u_00000005FA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[383*12+:12]), .o_data(C[127][1]), .i_clk(i_clk));
Mul0000000001  u_00000005FB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[639*12+:12]), .o_data(A[127][2]), .i_clk(i_clk));
Mul0000000001  u_00000005FC_Mul0000000001(.i_data_1(c_plus_d[127][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[127][2]), .i_clk(i_clk));
Mul0000000001  u_00000005FD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[639*12+:12]), .o_data(C[127][2]), .i_clk(i_clk));
Mul0000000001  u_00000005FE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[895*12+:12]), .o_data(A[127][3]), .i_clk(i_clk));
Mul0000000001  u_00000005FF_Mul0000000001(.i_data_1(c_plus_d[127][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[127][3]), .i_clk(i_clk));
Mul0000000001  u_0000000600_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[895*12+:12]), .o_data(C[127][3]), .i_clk(i_clk));
Mul0000000001  u_0000000601_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[128*12+:12]), .o_data(A[128][0]), .i_clk(i_clk));
Mul0000000001  u_0000000602_Mul0000000001(.i_data_1(c_plus_d[128][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[128][0]), .i_clk(i_clk));
Mul0000000001  u_0000000603_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[128*12+:12]), .o_data(C[128][0]), .i_clk(i_clk));
Mul0000000001  u_0000000604_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[384*12+:12]), .o_data(A[128][1]), .i_clk(i_clk));
Mul0000000001  u_0000000605_Mul0000000001(.i_data_1(c_plus_d[128][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[128][1]), .i_clk(i_clk));
Mul0000000001  u_0000000606_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[384*12+:12]), .o_data(C[128][1]), .i_clk(i_clk));
Mul0000000001  u_0000000607_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[640*12+:12]), .o_data(A[128][2]), .i_clk(i_clk));
Mul0000000001  u_0000000608_Mul0000000001(.i_data_1(c_plus_d[128][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[128][2]), .i_clk(i_clk));
Mul0000000001  u_0000000609_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[640*12+:12]), .o_data(C[128][2]), .i_clk(i_clk));
Mul0000000001  u_000000060A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[896*12+:12]), .o_data(A[128][3]), .i_clk(i_clk));
Mul0000000001  u_000000060B_Mul0000000001(.i_data_1(c_plus_d[128][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[128][3]), .i_clk(i_clk));
Mul0000000001  u_000000060C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[896*12+:12]), .o_data(C[128][3]), .i_clk(i_clk));
Mul0000000001  u_000000060D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[129*12+:12]), .o_data(A[129][0]), .i_clk(i_clk));
Mul0000000001  u_000000060E_Mul0000000001(.i_data_1(c_plus_d[129][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[129][0]), .i_clk(i_clk));
Mul0000000001  u_000000060F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[129*12+:12]), .o_data(C[129][0]), .i_clk(i_clk));
Mul0000000001  u_0000000610_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[385*12+:12]), .o_data(A[129][1]), .i_clk(i_clk));
Mul0000000001  u_0000000611_Mul0000000001(.i_data_1(c_plus_d[129][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[129][1]), .i_clk(i_clk));
Mul0000000001  u_0000000612_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[385*12+:12]), .o_data(C[129][1]), .i_clk(i_clk));
Mul0000000001  u_0000000613_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[641*12+:12]), .o_data(A[129][2]), .i_clk(i_clk));
Mul0000000001  u_0000000614_Mul0000000001(.i_data_1(c_plus_d[129][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[129][2]), .i_clk(i_clk));
Mul0000000001  u_0000000615_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[641*12+:12]), .o_data(C[129][2]), .i_clk(i_clk));
Mul0000000001  u_0000000616_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[897*12+:12]), .o_data(A[129][3]), .i_clk(i_clk));
Mul0000000001  u_0000000617_Mul0000000001(.i_data_1(c_plus_d[129][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[129][3]), .i_clk(i_clk));
Mul0000000001  u_0000000618_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[897*12+:12]), .o_data(C[129][3]), .i_clk(i_clk));
Mul0000000001  u_0000000619_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[130*12+:12]), .o_data(A[130][0]), .i_clk(i_clk));
Mul0000000001  u_000000061A_Mul0000000001(.i_data_1(c_plus_d[130][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[130][0]), .i_clk(i_clk));
Mul0000000001  u_000000061B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[130*12+:12]), .o_data(C[130][0]), .i_clk(i_clk));
Mul0000000001  u_000000061C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[386*12+:12]), .o_data(A[130][1]), .i_clk(i_clk));
Mul0000000001  u_000000061D_Mul0000000001(.i_data_1(c_plus_d[130][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[130][1]), .i_clk(i_clk));
Mul0000000001  u_000000061E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[386*12+:12]), .o_data(C[130][1]), .i_clk(i_clk));
Mul0000000001  u_000000061F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[642*12+:12]), .o_data(A[130][2]), .i_clk(i_clk));
Mul0000000001  u_0000000620_Mul0000000001(.i_data_1(c_plus_d[130][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[130][2]), .i_clk(i_clk));
Mul0000000001  u_0000000621_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[642*12+:12]), .o_data(C[130][2]), .i_clk(i_clk));
Mul0000000001  u_0000000622_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[898*12+:12]), .o_data(A[130][3]), .i_clk(i_clk));
Mul0000000001  u_0000000623_Mul0000000001(.i_data_1(c_plus_d[130][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[130][3]), .i_clk(i_clk));
Mul0000000001  u_0000000624_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[898*12+:12]), .o_data(C[130][3]), .i_clk(i_clk));
Mul0000000001  u_0000000625_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[131*12+:12]), .o_data(A[131][0]), .i_clk(i_clk));
Mul0000000001  u_0000000626_Mul0000000001(.i_data_1(c_plus_d[131][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[131][0]), .i_clk(i_clk));
Mul0000000001  u_0000000627_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[131*12+:12]), .o_data(C[131][0]), .i_clk(i_clk));
Mul0000000001  u_0000000628_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[387*12+:12]), .o_data(A[131][1]), .i_clk(i_clk));
Mul0000000001  u_0000000629_Mul0000000001(.i_data_1(c_plus_d[131][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[131][1]), .i_clk(i_clk));
Mul0000000001  u_000000062A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[387*12+:12]), .o_data(C[131][1]), .i_clk(i_clk));
Mul0000000001  u_000000062B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[643*12+:12]), .o_data(A[131][2]), .i_clk(i_clk));
Mul0000000001  u_000000062C_Mul0000000001(.i_data_1(c_plus_d[131][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[131][2]), .i_clk(i_clk));
Mul0000000001  u_000000062D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[643*12+:12]), .o_data(C[131][2]), .i_clk(i_clk));
Mul0000000001  u_000000062E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[899*12+:12]), .o_data(A[131][3]), .i_clk(i_clk));
Mul0000000001  u_000000062F_Mul0000000001(.i_data_1(c_plus_d[131][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[131][3]), .i_clk(i_clk));
Mul0000000001  u_0000000630_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[899*12+:12]), .o_data(C[131][3]), .i_clk(i_clk));
Mul0000000001  u_0000000631_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[132*12+:12]), .o_data(A[132][0]), .i_clk(i_clk));
Mul0000000001  u_0000000632_Mul0000000001(.i_data_1(c_plus_d[132][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[132][0]), .i_clk(i_clk));
Mul0000000001  u_0000000633_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[132*12+:12]), .o_data(C[132][0]), .i_clk(i_clk));
Mul0000000001  u_0000000634_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[388*12+:12]), .o_data(A[132][1]), .i_clk(i_clk));
Mul0000000001  u_0000000635_Mul0000000001(.i_data_1(c_plus_d[132][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[132][1]), .i_clk(i_clk));
Mul0000000001  u_0000000636_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[388*12+:12]), .o_data(C[132][1]), .i_clk(i_clk));
Mul0000000001  u_0000000637_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[644*12+:12]), .o_data(A[132][2]), .i_clk(i_clk));
Mul0000000001  u_0000000638_Mul0000000001(.i_data_1(c_plus_d[132][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[132][2]), .i_clk(i_clk));
Mul0000000001  u_0000000639_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[644*12+:12]), .o_data(C[132][2]), .i_clk(i_clk));
Mul0000000001  u_000000063A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[900*12+:12]), .o_data(A[132][3]), .i_clk(i_clk));
Mul0000000001  u_000000063B_Mul0000000001(.i_data_1(c_plus_d[132][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[132][3]), .i_clk(i_clk));
Mul0000000001  u_000000063C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[900*12+:12]), .o_data(C[132][3]), .i_clk(i_clk));
Mul0000000001  u_000000063D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[133*12+:12]), .o_data(A[133][0]), .i_clk(i_clk));
Mul0000000001  u_000000063E_Mul0000000001(.i_data_1(c_plus_d[133][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[133][0]), .i_clk(i_clk));
Mul0000000001  u_000000063F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[133*12+:12]), .o_data(C[133][0]), .i_clk(i_clk));
Mul0000000001  u_0000000640_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[389*12+:12]), .o_data(A[133][1]), .i_clk(i_clk));
Mul0000000001  u_0000000641_Mul0000000001(.i_data_1(c_plus_d[133][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[133][1]), .i_clk(i_clk));
Mul0000000001  u_0000000642_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[389*12+:12]), .o_data(C[133][1]), .i_clk(i_clk));
Mul0000000001  u_0000000643_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[645*12+:12]), .o_data(A[133][2]), .i_clk(i_clk));
Mul0000000001  u_0000000644_Mul0000000001(.i_data_1(c_plus_d[133][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[133][2]), .i_clk(i_clk));
Mul0000000001  u_0000000645_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[645*12+:12]), .o_data(C[133][2]), .i_clk(i_clk));
Mul0000000001  u_0000000646_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[901*12+:12]), .o_data(A[133][3]), .i_clk(i_clk));
Mul0000000001  u_0000000647_Mul0000000001(.i_data_1(c_plus_d[133][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[133][3]), .i_clk(i_clk));
Mul0000000001  u_0000000648_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[901*12+:12]), .o_data(C[133][3]), .i_clk(i_clk));
Mul0000000001  u_0000000649_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[134*12+:12]), .o_data(A[134][0]), .i_clk(i_clk));
Mul0000000001  u_000000064A_Mul0000000001(.i_data_1(c_plus_d[134][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[134][0]), .i_clk(i_clk));
Mul0000000001  u_000000064B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[134*12+:12]), .o_data(C[134][0]), .i_clk(i_clk));
Mul0000000001  u_000000064C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[390*12+:12]), .o_data(A[134][1]), .i_clk(i_clk));
Mul0000000001  u_000000064D_Mul0000000001(.i_data_1(c_plus_d[134][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[134][1]), .i_clk(i_clk));
Mul0000000001  u_000000064E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[390*12+:12]), .o_data(C[134][1]), .i_clk(i_clk));
Mul0000000001  u_000000064F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[646*12+:12]), .o_data(A[134][2]), .i_clk(i_clk));
Mul0000000001  u_0000000650_Mul0000000001(.i_data_1(c_plus_d[134][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[134][2]), .i_clk(i_clk));
Mul0000000001  u_0000000651_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[646*12+:12]), .o_data(C[134][2]), .i_clk(i_clk));
Mul0000000001  u_0000000652_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[902*12+:12]), .o_data(A[134][3]), .i_clk(i_clk));
Mul0000000001  u_0000000653_Mul0000000001(.i_data_1(c_plus_d[134][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[134][3]), .i_clk(i_clk));
Mul0000000001  u_0000000654_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[902*12+:12]), .o_data(C[134][3]), .i_clk(i_clk));
Mul0000000001  u_0000000655_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[135*12+:12]), .o_data(A[135][0]), .i_clk(i_clk));
Mul0000000001  u_0000000656_Mul0000000001(.i_data_1(c_plus_d[135][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[135][0]), .i_clk(i_clk));
Mul0000000001  u_0000000657_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[135*12+:12]), .o_data(C[135][0]), .i_clk(i_clk));
Mul0000000001  u_0000000658_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[391*12+:12]), .o_data(A[135][1]), .i_clk(i_clk));
Mul0000000001  u_0000000659_Mul0000000001(.i_data_1(c_plus_d[135][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[135][1]), .i_clk(i_clk));
Mul0000000001  u_000000065A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[391*12+:12]), .o_data(C[135][1]), .i_clk(i_clk));
Mul0000000001  u_000000065B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[647*12+:12]), .o_data(A[135][2]), .i_clk(i_clk));
Mul0000000001  u_000000065C_Mul0000000001(.i_data_1(c_plus_d[135][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[135][2]), .i_clk(i_clk));
Mul0000000001  u_000000065D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[647*12+:12]), .o_data(C[135][2]), .i_clk(i_clk));
Mul0000000001  u_000000065E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[903*12+:12]), .o_data(A[135][3]), .i_clk(i_clk));
Mul0000000001  u_000000065F_Mul0000000001(.i_data_1(c_plus_d[135][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[135][3]), .i_clk(i_clk));
Mul0000000001  u_0000000660_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[903*12+:12]), .o_data(C[135][3]), .i_clk(i_clk));
Mul0000000001  u_0000000661_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[136*12+:12]), .o_data(A[136][0]), .i_clk(i_clk));
Mul0000000001  u_0000000662_Mul0000000001(.i_data_1(c_plus_d[136][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[136][0]), .i_clk(i_clk));
Mul0000000001  u_0000000663_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[136*12+:12]), .o_data(C[136][0]), .i_clk(i_clk));
Mul0000000001  u_0000000664_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[392*12+:12]), .o_data(A[136][1]), .i_clk(i_clk));
Mul0000000001  u_0000000665_Mul0000000001(.i_data_1(c_plus_d[136][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[136][1]), .i_clk(i_clk));
Mul0000000001  u_0000000666_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[392*12+:12]), .o_data(C[136][1]), .i_clk(i_clk));
Mul0000000001  u_0000000667_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[648*12+:12]), .o_data(A[136][2]), .i_clk(i_clk));
Mul0000000001  u_0000000668_Mul0000000001(.i_data_1(c_plus_d[136][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[136][2]), .i_clk(i_clk));
Mul0000000001  u_0000000669_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[648*12+:12]), .o_data(C[136][2]), .i_clk(i_clk));
Mul0000000001  u_000000066A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[904*12+:12]), .o_data(A[136][3]), .i_clk(i_clk));
Mul0000000001  u_000000066B_Mul0000000001(.i_data_1(c_plus_d[136][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[136][3]), .i_clk(i_clk));
Mul0000000001  u_000000066C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[904*12+:12]), .o_data(C[136][3]), .i_clk(i_clk));
Mul0000000001  u_000000066D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[137*12+:12]), .o_data(A[137][0]), .i_clk(i_clk));
Mul0000000001  u_000000066E_Mul0000000001(.i_data_1(c_plus_d[137][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[137][0]), .i_clk(i_clk));
Mul0000000001  u_000000066F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[137*12+:12]), .o_data(C[137][0]), .i_clk(i_clk));
Mul0000000001  u_0000000670_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[393*12+:12]), .o_data(A[137][1]), .i_clk(i_clk));
Mul0000000001  u_0000000671_Mul0000000001(.i_data_1(c_plus_d[137][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[137][1]), .i_clk(i_clk));
Mul0000000001  u_0000000672_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[393*12+:12]), .o_data(C[137][1]), .i_clk(i_clk));
Mul0000000001  u_0000000673_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[649*12+:12]), .o_data(A[137][2]), .i_clk(i_clk));
Mul0000000001  u_0000000674_Mul0000000001(.i_data_1(c_plus_d[137][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[137][2]), .i_clk(i_clk));
Mul0000000001  u_0000000675_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[649*12+:12]), .o_data(C[137][2]), .i_clk(i_clk));
Mul0000000001  u_0000000676_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[905*12+:12]), .o_data(A[137][3]), .i_clk(i_clk));
Mul0000000001  u_0000000677_Mul0000000001(.i_data_1(c_plus_d[137][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[137][3]), .i_clk(i_clk));
Mul0000000001  u_0000000678_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[905*12+:12]), .o_data(C[137][3]), .i_clk(i_clk));
Mul0000000001  u_0000000679_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[138*12+:12]), .o_data(A[138][0]), .i_clk(i_clk));
Mul0000000001  u_000000067A_Mul0000000001(.i_data_1(c_plus_d[138][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[138][0]), .i_clk(i_clk));
Mul0000000001  u_000000067B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[138*12+:12]), .o_data(C[138][0]), .i_clk(i_clk));
Mul0000000001  u_000000067C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[394*12+:12]), .o_data(A[138][1]), .i_clk(i_clk));
Mul0000000001  u_000000067D_Mul0000000001(.i_data_1(c_plus_d[138][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[138][1]), .i_clk(i_clk));
Mul0000000001  u_000000067E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[394*12+:12]), .o_data(C[138][1]), .i_clk(i_clk));
Mul0000000001  u_000000067F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[650*12+:12]), .o_data(A[138][2]), .i_clk(i_clk));
Mul0000000001  u_0000000680_Mul0000000001(.i_data_1(c_plus_d[138][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[138][2]), .i_clk(i_clk));
Mul0000000001  u_0000000681_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[650*12+:12]), .o_data(C[138][2]), .i_clk(i_clk));
Mul0000000001  u_0000000682_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[906*12+:12]), .o_data(A[138][3]), .i_clk(i_clk));
Mul0000000001  u_0000000683_Mul0000000001(.i_data_1(c_plus_d[138][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[138][3]), .i_clk(i_clk));
Mul0000000001  u_0000000684_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[906*12+:12]), .o_data(C[138][3]), .i_clk(i_clk));
Mul0000000001  u_0000000685_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[139*12+:12]), .o_data(A[139][0]), .i_clk(i_clk));
Mul0000000001  u_0000000686_Mul0000000001(.i_data_1(c_plus_d[139][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[139][0]), .i_clk(i_clk));
Mul0000000001  u_0000000687_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[139*12+:12]), .o_data(C[139][0]), .i_clk(i_clk));
Mul0000000001  u_0000000688_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[395*12+:12]), .o_data(A[139][1]), .i_clk(i_clk));
Mul0000000001  u_0000000689_Mul0000000001(.i_data_1(c_plus_d[139][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[139][1]), .i_clk(i_clk));
Mul0000000001  u_000000068A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[395*12+:12]), .o_data(C[139][1]), .i_clk(i_clk));
Mul0000000001  u_000000068B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[651*12+:12]), .o_data(A[139][2]), .i_clk(i_clk));
Mul0000000001  u_000000068C_Mul0000000001(.i_data_1(c_plus_d[139][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[139][2]), .i_clk(i_clk));
Mul0000000001  u_000000068D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[651*12+:12]), .o_data(C[139][2]), .i_clk(i_clk));
Mul0000000001  u_000000068E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[907*12+:12]), .o_data(A[139][3]), .i_clk(i_clk));
Mul0000000001  u_000000068F_Mul0000000001(.i_data_1(c_plus_d[139][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[139][3]), .i_clk(i_clk));
Mul0000000001  u_0000000690_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[907*12+:12]), .o_data(C[139][3]), .i_clk(i_clk));
Mul0000000001  u_0000000691_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[140*12+:12]), .o_data(A[140][0]), .i_clk(i_clk));
Mul0000000001  u_0000000692_Mul0000000001(.i_data_1(c_plus_d[140][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[140][0]), .i_clk(i_clk));
Mul0000000001  u_0000000693_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[140*12+:12]), .o_data(C[140][0]), .i_clk(i_clk));
Mul0000000001  u_0000000694_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[396*12+:12]), .o_data(A[140][1]), .i_clk(i_clk));
Mul0000000001  u_0000000695_Mul0000000001(.i_data_1(c_plus_d[140][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[140][1]), .i_clk(i_clk));
Mul0000000001  u_0000000696_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[396*12+:12]), .o_data(C[140][1]), .i_clk(i_clk));
Mul0000000001  u_0000000697_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[652*12+:12]), .o_data(A[140][2]), .i_clk(i_clk));
Mul0000000001  u_0000000698_Mul0000000001(.i_data_1(c_plus_d[140][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[140][2]), .i_clk(i_clk));
Mul0000000001  u_0000000699_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[652*12+:12]), .o_data(C[140][2]), .i_clk(i_clk));
Mul0000000001  u_000000069A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[908*12+:12]), .o_data(A[140][3]), .i_clk(i_clk));
Mul0000000001  u_000000069B_Mul0000000001(.i_data_1(c_plus_d[140][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[140][3]), .i_clk(i_clk));
Mul0000000001  u_000000069C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[908*12+:12]), .o_data(C[140][3]), .i_clk(i_clk));
Mul0000000001  u_000000069D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[141*12+:12]), .o_data(A[141][0]), .i_clk(i_clk));
Mul0000000001  u_000000069E_Mul0000000001(.i_data_1(c_plus_d[141][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[141][0]), .i_clk(i_clk));
Mul0000000001  u_000000069F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[141*12+:12]), .o_data(C[141][0]), .i_clk(i_clk));
Mul0000000001  u_00000006A0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[397*12+:12]), .o_data(A[141][1]), .i_clk(i_clk));
Mul0000000001  u_00000006A1_Mul0000000001(.i_data_1(c_plus_d[141][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[141][1]), .i_clk(i_clk));
Mul0000000001  u_00000006A2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[397*12+:12]), .o_data(C[141][1]), .i_clk(i_clk));
Mul0000000001  u_00000006A3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[653*12+:12]), .o_data(A[141][2]), .i_clk(i_clk));
Mul0000000001  u_00000006A4_Mul0000000001(.i_data_1(c_plus_d[141][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[141][2]), .i_clk(i_clk));
Mul0000000001  u_00000006A5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[653*12+:12]), .o_data(C[141][2]), .i_clk(i_clk));
Mul0000000001  u_00000006A6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[909*12+:12]), .o_data(A[141][3]), .i_clk(i_clk));
Mul0000000001  u_00000006A7_Mul0000000001(.i_data_1(c_plus_d[141][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[141][3]), .i_clk(i_clk));
Mul0000000001  u_00000006A8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[909*12+:12]), .o_data(C[141][3]), .i_clk(i_clk));
Mul0000000001  u_00000006A9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[142*12+:12]), .o_data(A[142][0]), .i_clk(i_clk));
Mul0000000001  u_00000006AA_Mul0000000001(.i_data_1(c_plus_d[142][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[142][0]), .i_clk(i_clk));
Mul0000000001  u_00000006AB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[142*12+:12]), .o_data(C[142][0]), .i_clk(i_clk));
Mul0000000001  u_00000006AC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[398*12+:12]), .o_data(A[142][1]), .i_clk(i_clk));
Mul0000000001  u_00000006AD_Mul0000000001(.i_data_1(c_plus_d[142][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[142][1]), .i_clk(i_clk));
Mul0000000001  u_00000006AE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[398*12+:12]), .o_data(C[142][1]), .i_clk(i_clk));
Mul0000000001  u_00000006AF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[654*12+:12]), .o_data(A[142][2]), .i_clk(i_clk));
Mul0000000001  u_00000006B0_Mul0000000001(.i_data_1(c_plus_d[142][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[142][2]), .i_clk(i_clk));
Mul0000000001  u_00000006B1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[654*12+:12]), .o_data(C[142][2]), .i_clk(i_clk));
Mul0000000001  u_00000006B2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[910*12+:12]), .o_data(A[142][3]), .i_clk(i_clk));
Mul0000000001  u_00000006B3_Mul0000000001(.i_data_1(c_plus_d[142][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[142][3]), .i_clk(i_clk));
Mul0000000001  u_00000006B4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[910*12+:12]), .o_data(C[142][3]), .i_clk(i_clk));
Mul0000000001  u_00000006B5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[143*12+:12]), .o_data(A[143][0]), .i_clk(i_clk));
Mul0000000001  u_00000006B6_Mul0000000001(.i_data_1(c_plus_d[143][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[143][0]), .i_clk(i_clk));
Mul0000000001  u_00000006B7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[143*12+:12]), .o_data(C[143][0]), .i_clk(i_clk));
Mul0000000001  u_00000006B8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[399*12+:12]), .o_data(A[143][1]), .i_clk(i_clk));
Mul0000000001  u_00000006B9_Mul0000000001(.i_data_1(c_plus_d[143][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[143][1]), .i_clk(i_clk));
Mul0000000001  u_00000006BA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[399*12+:12]), .o_data(C[143][1]), .i_clk(i_clk));
Mul0000000001  u_00000006BB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[655*12+:12]), .o_data(A[143][2]), .i_clk(i_clk));
Mul0000000001  u_00000006BC_Mul0000000001(.i_data_1(c_plus_d[143][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[143][2]), .i_clk(i_clk));
Mul0000000001  u_00000006BD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[655*12+:12]), .o_data(C[143][2]), .i_clk(i_clk));
Mul0000000001  u_00000006BE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[911*12+:12]), .o_data(A[143][3]), .i_clk(i_clk));
Mul0000000001  u_00000006BF_Mul0000000001(.i_data_1(c_plus_d[143][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[143][3]), .i_clk(i_clk));
Mul0000000001  u_00000006C0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[911*12+:12]), .o_data(C[143][3]), .i_clk(i_clk));
Mul0000000001  u_00000006C1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[144*12+:12]), .o_data(A[144][0]), .i_clk(i_clk));
Mul0000000001  u_00000006C2_Mul0000000001(.i_data_1(c_plus_d[144][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[144][0]), .i_clk(i_clk));
Mul0000000001  u_00000006C3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[144*12+:12]), .o_data(C[144][0]), .i_clk(i_clk));
Mul0000000001  u_00000006C4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[400*12+:12]), .o_data(A[144][1]), .i_clk(i_clk));
Mul0000000001  u_00000006C5_Mul0000000001(.i_data_1(c_plus_d[144][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[144][1]), .i_clk(i_clk));
Mul0000000001  u_00000006C6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[400*12+:12]), .o_data(C[144][1]), .i_clk(i_clk));
Mul0000000001  u_00000006C7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[656*12+:12]), .o_data(A[144][2]), .i_clk(i_clk));
Mul0000000001  u_00000006C8_Mul0000000001(.i_data_1(c_plus_d[144][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[144][2]), .i_clk(i_clk));
Mul0000000001  u_00000006C9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[656*12+:12]), .o_data(C[144][2]), .i_clk(i_clk));
Mul0000000001  u_00000006CA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[912*12+:12]), .o_data(A[144][3]), .i_clk(i_clk));
Mul0000000001  u_00000006CB_Mul0000000001(.i_data_1(c_plus_d[144][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[144][3]), .i_clk(i_clk));
Mul0000000001  u_00000006CC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[912*12+:12]), .o_data(C[144][3]), .i_clk(i_clk));
Mul0000000001  u_00000006CD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[145*12+:12]), .o_data(A[145][0]), .i_clk(i_clk));
Mul0000000001  u_00000006CE_Mul0000000001(.i_data_1(c_plus_d[145][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[145][0]), .i_clk(i_clk));
Mul0000000001  u_00000006CF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[145*12+:12]), .o_data(C[145][0]), .i_clk(i_clk));
Mul0000000001  u_00000006D0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[401*12+:12]), .o_data(A[145][1]), .i_clk(i_clk));
Mul0000000001  u_00000006D1_Mul0000000001(.i_data_1(c_plus_d[145][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[145][1]), .i_clk(i_clk));
Mul0000000001  u_00000006D2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[401*12+:12]), .o_data(C[145][1]), .i_clk(i_clk));
Mul0000000001  u_00000006D3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[657*12+:12]), .o_data(A[145][2]), .i_clk(i_clk));
Mul0000000001  u_00000006D4_Mul0000000001(.i_data_1(c_plus_d[145][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[145][2]), .i_clk(i_clk));
Mul0000000001  u_00000006D5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[657*12+:12]), .o_data(C[145][2]), .i_clk(i_clk));
Mul0000000001  u_00000006D6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[913*12+:12]), .o_data(A[145][3]), .i_clk(i_clk));
Mul0000000001  u_00000006D7_Mul0000000001(.i_data_1(c_plus_d[145][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[145][3]), .i_clk(i_clk));
Mul0000000001  u_00000006D8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[913*12+:12]), .o_data(C[145][3]), .i_clk(i_clk));
Mul0000000001  u_00000006D9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[146*12+:12]), .o_data(A[146][0]), .i_clk(i_clk));
Mul0000000001  u_00000006DA_Mul0000000001(.i_data_1(c_plus_d[146][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[146][0]), .i_clk(i_clk));
Mul0000000001  u_00000006DB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[146*12+:12]), .o_data(C[146][0]), .i_clk(i_clk));
Mul0000000001  u_00000006DC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[402*12+:12]), .o_data(A[146][1]), .i_clk(i_clk));
Mul0000000001  u_00000006DD_Mul0000000001(.i_data_1(c_plus_d[146][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[146][1]), .i_clk(i_clk));
Mul0000000001  u_00000006DE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[402*12+:12]), .o_data(C[146][1]), .i_clk(i_clk));
Mul0000000001  u_00000006DF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[658*12+:12]), .o_data(A[146][2]), .i_clk(i_clk));
Mul0000000001  u_00000006E0_Mul0000000001(.i_data_1(c_plus_d[146][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[146][2]), .i_clk(i_clk));
Mul0000000001  u_00000006E1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[658*12+:12]), .o_data(C[146][2]), .i_clk(i_clk));
Mul0000000001  u_00000006E2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[914*12+:12]), .o_data(A[146][3]), .i_clk(i_clk));
Mul0000000001  u_00000006E3_Mul0000000001(.i_data_1(c_plus_d[146][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[146][3]), .i_clk(i_clk));
Mul0000000001  u_00000006E4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[914*12+:12]), .o_data(C[146][3]), .i_clk(i_clk));
Mul0000000001  u_00000006E5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[147*12+:12]), .o_data(A[147][0]), .i_clk(i_clk));
Mul0000000001  u_00000006E6_Mul0000000001(.i_data_1(c_plus_d[147][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[147][0]), .i_clk(i_clk));
Mul0000000001  u_00000006E7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[147*12+:12]), .o_data(C[147][0]), .i_clk(i_clk));
Mul0000000001  u_00000006E8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[403*12+:12]), .o_data(A[147][1]), .i_clk(i_clk));
Mul0000000001  u_00000006E9_Mul0000000001(.i_data_1(c_plus_d[147][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[147][1]), .i_clk(i_clk));
Mul0000000001  u_00000006EA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[403*12+:12]), .o_data(C[147][1]), .i_clk(i_clk));
Mul0000000001  u_00000006EB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[659*12+:12]), .o_data(A[147][2]), .i_clk(i_clk));
Mul0000000001  u_00000006EC_Mul0000000001(.i_data_1(c_plus_d[147][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[147][2]), .i_clk(i_clk));
Mul0000000001  u_00000006ED_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[659*12+:12]), .o_data(C[147][2]), .i_clk(i_clk));
Mul0000000001  u_00000006EE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[915*12+:12]), .o_data(A[147][3]), .i_clk(i_clk));
Mul0000000001  u_00000006EF_Mul0000000001(.i_data_1(c_plus_d[147][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[147][3]), .i_clk(i_clk));
Mul0000000001  u_00000006F0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[915*12+:12]), .o_data(C[147][3]), .i_clk(i_clk));
Mul0000000001  u_00000006F1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[148*12+:12]), .o_data(A[148][0]), .i_clk(i_clk));
Mul0000000001  u_00000006F2_Mul0000000001(.i_data_1(c_plus_d[148][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[148][0]), .i_clk(i_clk));
Mul0000000001  u_00000006F3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[148*12+:12]), .o_data(C[148][0]), .i_clk(i_clk));
Mul0000000001  u_00000006F4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[404*12+:12]), .o_data(A[148][1]), .i_clk(i_clk));
Mul0000000001  u_00000006F5_Mul0000000001(.i_data_1(c_plus_d[148][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[148][1]), .i_clk(i_clk));
Mul0000000001  u_00000006F6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[404*12+:12]), .o_data(C[148][1]), .i_clk(i_clk));
Mul0000000001  u_00000006F7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[660*12+:12]), .o_data(A[148][2]), .i_clk(i_clk));
Mul0000000001  u_00000006F8_Mul0000000001(.i_data_1(c_plus_d[148][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[148][2]), .i_clk(i_clk));
Mul0000000001  u_00000006F9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[660*12+:12]), .o_data(C[148][2]), .i_clk(i_clk));
Mul0000000001  u_00000006FA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[916*12+:12]), .o_data(A[148][3]), .i_clk(i_clk));
Mul0000000001  u_00000006FB_Mul0000000001(.i_data_1(c_plus_d[148][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[148][3]), .i_clk(i_clk));
Mul0000000001  u_00000006FC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[916*12+:12]), .o_data(C[148][3]), .i_clk(i_clk));
Mul0000000001  u_00000006FD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[149*12+:12]), .o_data(A[149][0]), .i_clk(i_clk));
Mul0000000001  u_00000006FE_Mul0000000001(.i_data_1(c_plus_d[149][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[149][0]), .i_clk(i_clk));
Mul0000000001  u_00000006FF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[149*12+:12]), .o_data(C[149][0]), .i_clk(i_clk));
Mul0000000001  u_0000000700_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[405*12+:12]), .o_data(A[149][1]), .i_clk(i_clk));
Mul0000000001  u_0000000701_Mul0000000001(.i_data_1(c_plus_d[149][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[149][1]), .i_clk(i_clk));
Mul0000000001  u_0000000702_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[405*12+:12]), .o_data(C[149][1]), .i_clk(i_clk));
Mul0000000001  u_0000000703_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[661*12+:12]), .o_data(A[149][2]), .i_clk(i_clk));
Mul0000000001  u_0000000704_Mul0000000001(.i_data_1(c_plus_d[149][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[149][2]), .i_clk(i_clk));
Mul0000000001  u_0000000705_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[661*12+:12]), .o_data(C[149][2]), .i_clk(i_clk));
Mul0000000001  u_0000000706_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[917*12+:12]), .o_data(A[149][3]), .i_clk(i_clk));
Mul0000000001  u_0000000707_Mul0000000001(.i_data_1(c_plus_d[149][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[149][3]), .i_clk(i_clk));
Mul0000000001  u_0000000708_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[917*12+:12]), .o_data(C[149][3]), .i_clk(i_clk));
Mul0000000001  u_0000000709_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[150*12+:12]), .o_data(A[150][0]), .i_clk(i_clk));
Mul0000000001  u_000000070A_Mul0000000001(.i_data_1(c_plus_d[150][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[150][0]), .i_clk(i_clk));
Mul0000000001  u_000000070B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[150*12+:12]), .o_data(C[150][0]), .i_clk(i_clk));
Mul0000000001  u_000000070C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[406*12+:12]), .o_data(A[150][1]), .i_clk(i_clk));
Mul0000000001  u_000000070D_Mul0000000001(.i_data_1(c_plus_d[150][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[150][1]), .i_clk(i_clk));
Mul0000000001  u_000000070E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[406*12+:12]), .o_data(C[150][1]), .i_clk(i_clk));
Mul0000000001  u_000000070F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[662*12+:12]), .o_data(A[150][2]), .i_clk(i_clk));
Mul0000000001  u_0000000710_Mul0000000001(.i_data_1(c_plus_d[150][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[150][2]), .i_clk(i_clk));
Mul0000000001  u_0000000711_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[662*12+:12]), .o_data(C[150][2]), .i_clk(i_clk));
Mul0000000001  u_0000000712_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[918*12+:12]), .o_data(A[150][3]), .i_clk(i_clk));
Mul0000000001  u_0000000713_Mul0000000001(.i_data_1(c_plus_d[150][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[150][3]), .i_clk(i_clk));
Mul0000000001  u_0000000714_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[918*12+:12]), .o_data(C[150][3]), .i_clk(i_clk));
Mul0000000001  u_0000000715_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[151*12+:12]), .o_data(A[151][0]), .i_clk(i_clk));
Mul0000000001  u_0000000716_Mul0000000001(.i_data_1(c_plus_d[151][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[151][0]), .i_clk(i_clk));
Mul0000000001  u_0000000717_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[151*12+:12]), .o_data(C[151][0]), .i_clk(i_clk));
Mul0000000001  u_0000000718_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[407*12+:12]), .o_data(A[151][1]), .i_clk(i_clk));
Mul0000000001  u_0000000719_Mul0000000001(.i_data_1(c_plus_d[151][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[151][1]), .i_clk(i_clk));
Mul0000000001  u_000000071A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[407*12+:12]), .o_data(C[151][1]), .i_clk(i_clk));
Mul0000000001  u_000000071B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[663*12+:12]), .o_data(A[151][2]), .i_clk(i_clk));
Mul0000000001  u_000000071C_Mul0000000001(.i_data_1(c_plus_d[151][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[151][2]), .i_clk(i_clk));
Mul0000000001  u_000000071D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[663*12+:12]), .o_data(C[151][2]), .i_clk(i_clk));
Mul0000000001  u_000000071E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[919*12+:12]), .o_data(A[151][3]), .i_clk(i_clk));
Mul0000000001  u_000000071F_Mul0000000001(.i_data_1(c_plus_d[151][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[151][3]), .i_clk(i_clk));
Mul0000000001  u_0000000720_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[919*12+:12]), .o_data(C[151][3]), .i_clk(i_clk));
Mul0000000001  u_0000000721_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[152*12+:12]), .o_data(A[152][0]), .i_clk(i_clk));
Mul0000000001  u_0000000722_Mul0000000001(.i_data_1(c_plus_d[152][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[152][0]), .i_clk(i_clk));
Mul0000000001  u_0000000723_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[152*12+:12]), .o_data(C[152][0]), .i_clk(i_clk));
Mul0000000001  u_0000000724_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[408*12+:12]), .o_data(A[152][1]), .i_clk(i_clk));
Mul0000000001  u_0000000725_Mul0000000001(.i_data_1(c_plus_d[152][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[152][1]), .i_clk(i_clk));
Mul0000000001  u_0000000726_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[408*12+:12]), .o_data(C[152][1]), .i_clk(i_clk));
Mul0000000001  u_0000000727_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[664*12+:12]), .o_data(A[152][2]), .i_clk(i_clk));
Mul0000000001  u_0000000728_Mul0000000001(.i_data_1(c_plus_d[152][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[152][2]), .i_clk(i_clk));
Mul0000000001  u_0000000729_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[664*12+:12]), .o_data(C[152][2]), .i_clk(i_clk));
Mul0000000001  u_000000072A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[920*12+:12]), .o_data(A[152][3]), .i_clk(i_clk));
Mul0000000001  u_000000072B_Mul0000000001(.i_data_1(c_plus_d[152][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[152][3]), .i_clk(i_clk));
Mul0000000001  u_000000072C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[920*12+:12]), .o_data(C[152][3]), .i_clk(i_clk));
Mul0000000001  u_000000072D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[153*12+:12]), .o_data(A[153][0]), .i_clk(i_clk));
Mul0000000001  u_000000072E_Mul0000000001(.i_data_1(c_plus_d[153][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[153][0]), .i_clk(i_clk));
Mul0000000001  u_000000072F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[153*12+:12]), .o_data(C[153][0]), .i_clk(i_clk));
Mul0000000001  u_0000000730_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[409*12+:12]), .o_data(A[153][1]), .i_clk(i_clk));
Mul0000000001  u_0000000731_Mul0000000001(.i_data_1(c_plus_d[153][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[153][1]), .i_clk(i_clk));
Mul0000000001  u_0000000732_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[409*12+:12]), .o_data(C[153][1]), .i_clk(i_clk));
Mul0000000001  u_0000000733_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[665*12+:12]), .o_data(A[153][2]), .i_clk(i_clk));
Mul0000000001  u_0000000734_Mul0000000001(.i_data_1(c_plus_d[153][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[153][2]), .i_clk(i_clk));
Mul0000000001  u_0000000735_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[665*12+:12]), .o_data(C[153][2]), .i_clk(i_clk));
Mul0000000001  u_0000000736_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[921*12+:12]), .o_data(A[153][3]), .i_clk(i_clk));
Mul0000000001  u_0000000737_Mul0000000001(.i_data_1(c_plus_d[153][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[153][3]), .i_clk(i_clk));
Mul0000000001  u_0000000738_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[921*12+:12]), .o_data(C[153][3]), .i_clk(i_clk));
Mul0000000001  u_0000000739_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[154*12+:12]), .o_data(A[154][0]), .i_clk(i_clk));
Mul0000000001  u_000000073A_Mul0000000001(.i_data_1(c_plus_d[154][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[154][0]), .i_clk(i_clk));
Mul0000000001  u_000000073B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[154*12+:12]), .o_data(C[154][0]), .i_clk(i_clk));
Mul0000000001  u_000000073C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[410*12+:12]), .o_data(A[154][1]), .i_clk(i_clk));
Mul0000000001  u_000000073D_Mul0000000001(.i_data_1(c_plus_d[154][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[154][1]), .i_clk(i_clk));
Mul0000000001  u_000000073E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[410*12+:12]), .o_data(C[154][1]), .i_clk(i_clk));
Mul0000000001  u_000000073F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[666*12+:12]), .o_data(A[154][2]), .i_clk(i_clk));
Mul0000000001  u_0000000740_Mul0000000001(.i_data_1(c_plus_d[154][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[154][2]), .i_clk(i_clk));
Mul0000000001  u_0000000741_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[666*12+:12]), .o_data(C[154][2]), .i_clk(i_clk));
Mul0000000001  u_0000000742_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[922*12+:12]), .o_data(A[154][3]), .i_clk(i_clk));
Mul0000000001  u_0000000743_Mul0000000001(.i_data_1(c_plus_d[154][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[154][3]), .i_clk(i_clk));
Mul0000000001  u_0000000744_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[922*12+:12]), .o_data(C[154][3]), .i_clk(i_clk));
Mul0000000001  u_0000000745_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[155*12+:12]), .o_data(A[155][0]), .i_clk(i_clk));
Mul0000000001  u_0000000746_Mul0000000001(.i_data_1(c_plus_d[155][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[155][0]), .i_clk(i_clk));
Mul0000000001  u_0000000747_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[155*12+:12]), .o_data(C[155][0]), .i_clk(i_clk));
Mul0000000001  u_0000000748_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[411*12+:12]), .o_data(A[155][1]), .i_clk(i_clk));
Mul0000000001  u_0000000749_Mul0000000001(.i_data_1(c_plus_d[155][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[155][1]), .i_clk(i_clk));
Mul0000000001  u_000000074A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[411*12+:12]), .o_data(C[155][1]), .i_clk(i_clk));
Mul0000000001  u_000000074B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[667*12+:12]), .o_data(A[155][2]), .i_clk(i_clk));
Mul0000000001  u_000000074C_Mul0000000001(.i_data_1(c_plus_d[155][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[155][2]), .i_clk(i_clk));
Mul0000000001  u_000000074D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[667*12+:12]), .o_data(C[155][2]), .i_clk(i_clk));
Mul0000000001  u_000000074E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[923*12+:12]), .o_data(A[155][3]), .i_clk(i_clk));
Mul0000000001  u_000000074F_Mul0000000001(.i_data_1(c_plus_d[155][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[155][3]), .i_clk(i_clk));
Mul0000000001  u_0000000750_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[923*12+:12]), .o_data(C[155][3]), .i_clk(i_clk));
Mul0000000001  u_0000000751_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[156*12+:12]), .o_data(A[156][0]), .i_clk(i_clk));
Mul0000000001  u_0000000752_Mul0000000001(.i_data_1(c_plus_d[156][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[156][0]), .i_clk(i_clk));
Mul0000000001  u_0000000753_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[156*12+:12]), .o_data(C[156][0]), .i_clk(i_clk));
Mul0000000001  u_0000000754_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[412*12+:12]), .o_data(A[156][1]), .i_clk(i_clk));
Mul0000000001  u_0000000755_Mul0000000001(.i_data_1(c_plus_d[156][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[156][1]), .i_clk(i_clk));
Mul0000000001  u_0000000756_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[412*12+:12]), .o_data(C[156][1]), .i_clk(i_clk));
Mul0000000001  u_0000000757_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[668*12+:12]), .o_data(A[156][2]), .i_clk(i_clk));
Mul0000000001  u_0000000758_Mul0000000001(.i_data_1(c_plus_d[156][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[156][2]), .i_clk(i_clk));
Mul0000000001  u_0000000759_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[668*12+:12]), .o_data(C[156][2]), .i_clk(i_clk));
Mul0000000001  u_000000075A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[924*12+:12]), .o_data(A[156][3]), .i_clk(i_clk));
Mul0000000001  u_000000075B_Mul0000000001(.i_data_1(c_plus_d[156][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[156][3]), .i_clk(i_clk));
Mul0000000001  u_000000075C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[924*12+:12]), .o_data(C[156][3]), .i_clk(i_clk));
Mul0000000001  u_000000075D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[157*12+:12]), .o_data(A[157][0]), .i_clk(i_clk));
Mul0000000001  u_000000075E_Mul0000000001(.i_data_1(c_plus_d[157][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[157][0]), .i_clk(i_clk));
Mul0000000001  u_000000075F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[157*12+:12]), .o_data(C[157][0]), .i_clk(i_clk));
Mul0000000001  u_0000000760_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[413*12+:12]), .o_data(A[157][1]), .i_clk(i_clk));
Mul0000000001  u_0000000761_Mul0000000001(.i_data_1(c_plus_d[157][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[157][1]), .i_clk(i_clk));
Mul0000000001  u_0000000762_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[413*12+:12]), .o_data(C[157][1]), .i_clk(i_clk));
Mul0000000001  u_0000000763_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[669*12+:12]), .o_data(A[157][2]), .i_clk(i_clk));
Mul0000000001  u_0000000764_Mul0000000001(.i_data_1(c_plus_d[157][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[157][2]), .i_clk(i_clk));
Mul0000000001  u_0000000765_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[669*12+:12]), .o_data(C[157][2]), .i_clk(i_clk));
Mul0000000001  u_0000000766_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[925*12+:12]), .o_data(A[157][3]), .i_clk(i_clk));
Mul0000000001  u_0000000767_Mul0000000001(.i_data_1(c_plus_d[157][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[157][3]), .i_clk(i_clk));
Mul0000000001  u_0000000768_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[925*12+:12]), .o_data(C[157][3]), .i_clk(i_clk));
Mul0000000001  u_0000000769_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[158*12+:12]), .o_data(A[158][0]), .i_clk(i_clk));
Mul0000000001  u_000000076A_Mul0000000001(.i_data_1(c_plus_d[158][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[158][0]), .i_clk(i_clk));
Mul0000000001  u_000000076B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[158*12+:12]), .o_data(C[158][0]), .i_clk(i_clk));
Mul0000000001  u_000000076C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[414*12+:12]), .o_data(A[158][1]), .i_clk(i_clk));
Mul0000000001  u_000000076D_Mul0000000001(.i_data_1(c_plus_d[158][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[158][1]), .i_clk(i_clk));
Mul0000000001  u_000000076E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[414*12+:12]), .o_data(C[158][1]), .i_clk(i_clk));
Mul0000000001  u_000000076F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[670*12+:12]), .o_data(A[158][2]), .i_clk(i_clk));
Mul0000000001  u_0000000770_Mul0000000001(.i_data_1(c_plus_d[158][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[158][2]), .i_clk(i_clk));
Mul0000000001  u_0000000771_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[670*12+:12]), .o_data(C[158][2]), .i_clk(i_clk));
Mul0000000001  u_0000000772_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[926*12+:12]), .o_data(A[158][3]), .i_clk(i_clk));
Mul0000000001  u_0000000773_Mul0000000001(.i_data_1(c_plus_d[158][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[158][3]), .i_clk(i_clk));
Mul0000000001  u_0000000774_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[926*12+:12]), .o_data(C[158][3]), .i_clk(i_clk));
Mul0000000001  u_0000000775_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[159*12+:12]), .o_data(A[159][0]), .i_clk(i_clk));
Mul0000000001  u_0000000776_Mul0000000001(.i_data_1(c_plus_d[159][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[159][0]), .i_clk(i_clk));
Mul0000000001  u_0000000777_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[159*12+:12]), .o_data(C[159][0]), .i_clk(i_clk));
Mul0000000001  u_0000000778_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[415*12+:12]), .o_data(A[159][1]), .i_clk(i_clk));
Mul0000000001  u_0000000779_Mul0000000001(.i_data_1(c_plus_d[159][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[159][1]), .i_clk(i_clk));
Mul0000000001  u_000000077A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[415*12+:12]), .o_data(C[159][1]), .i_clk(i_clk));
Mul0000000001  u_000000077B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[671*12+:12]), .o_data(A[159][2]), .i_clk(i_clk));
Mul0000000001  u_000000077C_Mul0000000001(.i_data_1(c_plus_d[159][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[159][2]), .i_clk(i_clk));
Mul0000000001  u_000000077D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[671*12+:12]), .o_data(C[159][2]), .i_clk(i_clk));
Mul0000000001  u_000000077E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[927*12+:12]), .o_data(A[159][3]), .i_clk(i_clk));
Mul0000000001  u_000000077F_Mul0000000001(.i_data_1(c_plus_d[159][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[159][3]), .i_clk(i_clk));
Mul0000000001  u_0000000780_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[927*12+:12]), .o_data(C[159][3]), .i_clk(i_clk));
Mul0000000001  u_0000000781_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[160*12+:12]), .o_data(A[160][0]), .i_clk(i_clk));
Mul0000000001  u_0000000782_Mul0000000001(.i_data_1(c_plus_d[160][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[160][0]), .i_clk(i_clk));
Mul0000000001  u_0000000783_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[160*12+:12]), .o_data(C[160][0]), .i_clk(i_clk));
Mul0000000001  u_0000000784_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[416*12+:12]), .o_data(A[160][1]), .i_clk(i_clk));
Mul0000000001  u_0000000785_Mul0000000001(.i_data_1(c_plus_d[160][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[160][1]), .i_clk(i_clk));
Mul0000000001  u_0000000786_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[416*12+:12]), .o_data(C[160][1]), .i_clk(i_clk));
Mul0000000001  u_0000000787_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[672*12+:12]), .o_data(A[160][2]), .i_clk(i_clk));
Mul0000000001  u_0000000788_Mul0000000001(.i_data_1(c_plus_d[160][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[160][2]), .i_clk(i_clk));
Mul0000000001  u_0000000789_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[672*12+:12]), .o_data(C[160][2]), .i_clk(i_clk));
Mul0000000001  u_000000078A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[928*12+:12]), .o_data(A[160][3]), .i_clk(i_clk));
Mul0000000001  u_000000078B_Mul0000000001(.i_data_1(c_plus_d[160][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[160][3]), .i_clk(i_clk));
Mul0000000001  u_000000078C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[928*12+:12]), .o_data(C[160][3]), .i_clk(i_clk));
Mul0000000001  u_000000078D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[161*12+:12]), .o_data(A[161][0]), .i_clk(i_clk));
Mul0000000001  u_000000078E_Mul0000000001(.i_data_1(c_plus_d[161][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[161][0]), .i_clk(i_clk));
Mul0000000001  u_000000078F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[161*12+:12]), .o_data(C[161][0]), .i_clk(i_clk));
Mul0000000001  u_0000000790_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[417*12+:12]), .o_data(A[161][1]), .i_clk(i_clk));
Mul0000000001  u_0000000791_Mul0000000001(.i_data_1(c_plus_d[161][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[161][1]), .i_clk(i_clk));
Mul0000000001  u_0000000792_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[417*12+:12]), .o_data(C[161][1]), .i_clk(i_clk));
Mul0000000001  u_0000000793_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[673*12+:12]), .o_data(A[161][2]), .i_clk(i_clk));
Mul0000000001  u_0000000794_Mul0000000001(.i_data_1(c_plus_d[161][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[161][2]), .i_clk(i_clk));
Mul0000000001  u_0000000795_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[673*12+:12]), .o_data(C[161][2]), .i_clk(i_clk));
Mul0000000001  u_0000000796_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[929*12+:12]), .o_data(A[161][3]), .i_clk(i_clk));
Mul0000000001  u_0000000797_Mul0000000001(.i_data_1(c_plus_d[161][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[161][3]), .i_clk(i_clk));
Mul0000000001  u_0000000798_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[929*12+:12]), .o_data(C[161][3]), .i_clk(i_clk));
Mul0000000001  u_0000000799_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[162*12+:12]), .o_data(A[162][0]), .i_clk(i_clk));
Mul0000000001  u_000000079A_Mul0000000001(.i_data_1(c_plus_d[162][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[162][0]), .i_clk(i_clk));
Mul0000000001  u_000000079B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[162*12+:12]), .o_data(C[162][0]), .i_clk(i_clk));
Mul0000000001  u_000000079C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[418*12+:12]), .o_data(A[162][1]), .i_clk(i_clk));
Mul0000000001  u_000000079D_Mul0000000001(.i_data_1(c_plus_d[162][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[162][1]), .i_clk(i_clk));
Mul0000000001  u_000000079E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[418*12+:12]), .o_data(C[162][1]), .i_clk(i_clk));
Mul0000000001  u_000000079F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[674*12+:12]), .o_data(A[162][2]), .i_clk(i_clk));
Mul0000000001  u_00000007A0_Mul0000000001(.i_data_1(c_plus_d[162][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[162][2]), .i_clk(i_clk));
Mul0000000001  u_00000007A1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[674*12+:12]), .o_data(C[162][2]), .i_clk(i_clk));
Mul0000000001  u_00000007A2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[930*12+:12]), .o_data(A[162][3]), .i_clk(i_clk));
Mul0000000001  u_00000007A3_Mul0000000001(.i_data_1(c_plus_d[162][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[162][3]), .i_clk(i_clk));
Mul0000000001  u_00000007A4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[930*12+:12]), .o_data(C[162][3]), .i_clk(i_clk));
Mul0000000001  u_00000007A5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[163*12+:12]), .o_data(A[163][0]), .i_clk(i_clk));
Mul0000000001  u_00000007A6_Mul0000000001(.i_data_1(c_plus_d[163][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[163][0]), .i_clk(i_clk));
Mul0000000001  u_00000007A7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[163*12+:12]), .o_data(C[163][0]), .i_clk(i_clk));
Mul0000000001  u_00000007A8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[419*12+:12]), .o_data(A[163][1]), .i_clk(i_clk));
Mul0000000001  u_00000007A9_Mul0000000001(.i_data_1(c_plus_d[163][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[163][1]), .i_clk(i_clk));
Mul0000000001  u_00000007AA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[419*12+:12]), .o_data(C[163][1]), .i_clk(i_clk));
Mul0000000001  u_00000007AB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[675*12+:12]), .o_data(A[163][2]), .i_clk(i_clk));
Mul0000000001  u_00000007AC_Mul0000000001(.i_data_1(c_plus_d[163][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[163][2]), .i_clk(i_clk));
Mul0000000001  u_00000007AD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[675*12+:12]), .o_data(C[163][2]), .i_clk(i_clk));
Mul0000000001  u_00000007AE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[931*12+:12]), .o_data(A[163][3]), .i_clk(i_clk));
Mul0000000001  u_00000007AF_Mul0000000001(.i_data_1(c_plus_d[163][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[163][3]), .i_clk(i_clk));
Mul0000000001  u_00000007B0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[931*12+:12]), .o_data(C[163][3]), .i_clk(i_clk));
Mul0000000001  u_00000007B1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[164*12+:12]), .o_data(A[164][0]), .i_clk(i_clk));
Mul0000000001  u_00000007B2_Mul0000000001(.i_data_1(c_plus_d[164][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[164][0]), .i_clk(i_clk));
Mul0000000001  u_00000007B3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[164*12+:12]), .o_data(C[164][0]), .i_clk(i_clk));
Mul0000000001  u_00000007B4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[420*12+:12]), .o_data(A[164][1]), .i_clk(i_clk));
Mul0000000001  u_00000007B5_Mul0000000001(.i_data_1(c_plus_d[164][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[164][1]), .i_clk(i_clk));
Mul0000000001  u_00000007B6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[420*12+:12]), .o_data(C[164][1]), .i_clk(i_clk));
Mul0000000001  u_00000007B7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[676*12+:12]), .o_data(A[164][2]), .i_clk(i_clk));
Mul0000000001  u_00000007B8_Mul0000000001(.i_data_1(c_plus_d[164][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[164][2]), .i_clk(i_clk));
Mul0000000001  u_00000007B9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[676*12+:12]), .o_data(C[164][2]), .i_clk(i_clk));
Mul0000000001  u_00000007BA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[932*12+:12]), .o_data(A[164][3]), .i_clk(i_clk));
Mul0000000001  u_00000007BB_Mul0000000001(.i_data_1(c_plus_d[164][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[164][3]), .i_clk(i_clk));
Mul0000000001  u_00000007BC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[932*12+:12]), .o_data(C[164][3]), .i_clk(i_clk));
Mul0000000001  u_00000007BD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[165*12+:12]), .o_data(A[165][0]), .i_clk(i_clk));
Mul0000000001  u_00000007BE_Mul0000000001(.i_data_1(c_plus_d[165][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[165][0]), .i_clk(i_clk));
Mul0000000001  u_00000007BF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[165*12+:12]), .o_data(C[165][0]), .i_clk(i_clk));
Mul0000000001  u_00000007C0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[421*12+:12]), .o_data(A[165][1]), .i_clk(i_clk));
Mul0000000001  u_00000007C1_Mul0000000001(.i_data_1(c_plus_d[165][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[165][1]), .i_clk(i_clk));
Mul0000000001  u_00000007C2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[421*12+:12]), .o_data(C[165][1]), .i_clk(i_clk));
Mul0000000001  u_00000007C3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[677*12+:12]), .o_data(A[165][2]), .i_clk(i_clk));
Mul0000000001  u_00000007C4_Mul0000000001(.i_data_1(c_plus_d[165][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[165][2]), .i_clk(i_clk));
Mul0000000001  u_00000007C5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[677*12+:12]), .o_data(C[165][2]), .i_clk(i_clk));
Mul0000000001  u_00000007C6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[933*12+:12]), .o_data(A[165][3]), .i_clk(i_clk));
Mul0000000001  u_00000007C7_Mul0000000001(.i_data_1(c_plus_d[165][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[165][3]), .i_clk(i_clk));
Mul0000000001  u_00000007C8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[933*12+:12]), .o_data(C[165][3]), .i_clk(i_clk));
Mul0000000001  u_00000007C9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[166*12+:12]), .o_data(A[166][0]), .i_clk(i_clk));
Mul0000000001  u_00000007CA_Mul0000000001(.i_data_1(c_plus_d[166][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[166][0]), .i_clk(i_clk));
Mul0000000001  u_00000007CB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[166*12+:12]), .o_data(C[166][0]), .i_clk(i_clk));
Mul0000000001  u_00000007CC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[422*12+:12]), .o_data(A[166][1]), .i_clk(i_clk));
Mul0000000001  u_00000007CD_Mul0000000001(.i_data_1(c_plus_d[166][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[166][1]), .i_clk(i_clk));
Mul0000000001  u_00000007CE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[422*12+:12]), .o_data(C[166][1]), .i_clk(i_clk));
Mul0000000001  u_00000007CF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[678*12+:12]), .o_data(A[166][2]), .i_clk(i_clk));
Mul0000000001  u_00000007D0_Mul0000000001(.i_data_1(c_plus_d[166][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[166][2]), .i_clk(i_clk));
Mul0000000001  u_00000007D1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[678*12+:12]), .o_data(C[166][2]), .i_clk(i_clk));
Mul0000000001  u_00000007D2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[934*12+:12]), .o_data(A[166][3]), .i_clk(i_clk));
Mul0000000001  u_00000007D3_Mul0000000001(.i_data_1(c_plus_d[166][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[166][3]), .i_clk(i_clk));
Mul0000000001  u_00000007D4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[934*12+:12]), .o_data(C[166][3]), .i_clk(i_clk));
Mul0000000001  u_00000007D5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[167*12+:12]), .o_data(A[167][0]), .i_clk(i_clk));
Mul0000000001  u_00000007D6_Mul0000000001(.i_data_1(c_plus_d[167][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[167][0]), .i_clk(i_clk));
Mul0000000001  u_00000007D7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[167*12+:12]), .o_data(C[167][0]), .i_clk(i_clk));
Mul0000000001  u_00000007D8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[423*12+:12]), .o_data(A[167][1]), .i_clk(i_clk));
Mul0000000001  u_00000007D9_Mul0000000001(.i_data_1(c_plus_d[167][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[167][1]), .i_clk(i_clk));
Mul0000000001  u_00000007DA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[423*12+:12]), .o_data(C[167][1]), .i_clk(i_clk));
Mul0000000001  u_00000007DB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[679*12+:12]), .o_data(A[167][2]), .i_clk(i_clk));
Mul0000000001  u_00000007DC_Mul0000000001(.i_data_1(c_plus_d[167][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[167][2]), .i_clk(i_clk));
Mul0000000001  u_00000007DD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[679*12+:12]), .o_data(C[167][2]), .i_clk(i_clk));
Mul0000000001  u_00000007DE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[935*12+:12]), .o_data(A[167][3]), .i_clk(i_clk));
Mul0000000001  u_00000007DF_Mul0000000001(.i_data_1(c_plus_d[167][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[167][3]), .i_clk(i_clk));
Mul0000000001  u_00000007E0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[935*12+:12]), .o_data(C[167][3]), .i_clk(i_clk));
Mul0000000001  u_00000007E1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[168*12+:12]), .o_data(A[168][0]), .i_clk(i_clk));
Mul0000000001  u_00000007E2_Mul0000000001(.i_data_1(c_plus_d[168][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[168][0]), .i_clk(i_clk));
Mul0000000001  u_00000007E3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[168*12+:12]), .o_data(C[168][0]), .i_clk(i_clk));
Mul0000000001  u_00000007E4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[424*12+:12]), .o_data(A[168][1]), .i_clk(i_clk));
Mul0000000001  u_00000007E5_Mul0000000001(.i_data_1(c_plus_d[168][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[168][1]), .i_clk(i_clk));
Mul0000000001  u_00000007E6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[424*12+:12]), .o_data(C[168][1]), .i_clk(i_clk));
Mul0000000001  u_00000007E7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[680*12+:12]), .o_data(A[168][2]), .i_clk(i_clk));
Mul0000000001  u_00000007E8_Mul0000000001(.i_data_1(c_plus_d[168][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[168][2]), .i_clk(i_clk));
Mul0000000001  u_00000007E9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[680*12+:12]), .o_data(C[168][2]), .i_clk(i_clk));
Mul0000000001  u_00000007EA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[936*12+:12]), .o_data(A[168][3]), .i_clk(i_clk));
Mul0000000001  u_00000007EB_Mul0000000001(.i_data_1(c_plus_d[168][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[168][3]), .i_clk(i_clk));
Mul0000000001  u_00000007EC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[936*12+:12]), .o_data(C[168][3]), .i_clk(i_clk));
Mul0000000001  u_00000007ED_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[169*12+:12]), .o_data(A[169][0]), .i_clk(i_clk));
Mul0000000001  u_00000007EE_Mul0000000001(.i_data_1(c_plus_d[169][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[169][0]), .i_clk(i_clk));
Mul0000000001  u_00000007EF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[169*12+:12]), .o_data(C[169][0]), .i_clk(i_clk));
Mul0000000001  u_00000007F0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[425*12+:12]), .o_data(A[169][1]), .i_clk(i_clk));
Mul0000000001  u_00000007F1_Mul0000000001(.i_data_1(c_plus_d[169][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[169][1]), .i_clk(i_clk));
Mul0000000001  u_00000007F2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[425*12+:12]), .o_data(C[169][1]), .i_clk(i_clk));
Mul0000000001  u_00000007F3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[681*12+:12]), .o_data(A[169][2]), .i_clk(i_clk));
Mul0000000001  u_00000007F4_Mul0000000001(.i_data_1(c_plus_d[169][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[169][2]), .i_clk(i_clk));
Mul0000000001  u_00000007F5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[681*12+:12]), .o_data(C[169][2]), .i_clk(i_clk));
Mul0000000001  u_00000007F6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[937*12+:12]), .o_data(A[169][3]), .i_clk(i_clk));
Mul0000000001  u_00000007F7_Mul0000000001(.i_data_1(c_plus_d[169][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[169][3]), .i_clk(i_clk));
Mul0000000001  u_00000007F8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[937*12+:12]), .o_data(C[169][3]), .i_clk(i_clk));
Mul0000000001  u_00000007F9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[170*12+:12]), .o_data(A[170][0]), .i_clk(i_clk));
Mul0000000001  u_00000007FA_Mul0000000001(.i_data_1(c_plus_d[170][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[170][0]), .i_clk(i_clk));
Mul0000000001  u_00000007FB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[170*12+:12]), .o_data(C[170][0]), .i_clk(i_clk));
Mul0000000001  u_00000007FC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[426*12+:12]), .o_data(A[170][1]), .i_clk(i_clk));
Mul0000000001  u_00000007FD_Mul0000000001(.i_data_1(c_plus_d[170][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[170][1]), .i_clk(i_clk));
Mul0000000001  u_00000007FE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[426*12+:12]), .o_data(C[170][1]), .i_clk(i_clk));
Mul0000000001  u_00000007FF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[682*12+:12]), .o_data(A[170][2]), .i_clk(i_clk));
Mul0000000001  u_0000000800_Mul0000000001(.i_data_1(c_plus_d[170][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[170][2]), .i_clk(i_clk));
Mul0000000001  u_0000000801_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[682*12+:12]), .o_data(C[170][2]), .i_clk(i_clk));
Mul0000000001  u_0000000802_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[938*12+:12]), .o_data(A[170][3]), .i_clk(i_clk));
Mul0000000001  u_0000000803_Mul0000000001(.i_data_1(c_plus_d[170][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[170][3]), .i_clk(i_clk));
Mul0000000001  u_0000000804_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[938*12+:12]), .o_data(C[170][3]), .i_clk(i_clk));
Mul0000000001  u_0000000805_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[171*12+:12]), .o_data(A[171][0]), .i_clk(i_clk));
Mul0000000001  u_0000000806_Mul0000000001(.i_data_1(c_plus_d[171][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[171][0]), .i_clk(i_clk));
Mul0000000001  u_0000000807_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[171*12+:12]), .o_data(C[171][0]), .i_clk(i_clk));
Mul0000000001  u_0000000808_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[427*12+:12]), .o_data(A[171][1]), .i_clk(i_clk));
Mul0000000001  u_0000000809_Mul0000000001(.i_data_1(c_plus_d[171][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[171][1]), .i_clk(i_clk));
Mul0000000001  u_000000080A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[427*12+:12]), .o_data(C[171][1]), .i_clk(i_clk));
Mul0000000001  u_000000080B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[683*12+:12]), .o_data(A[171][2]), .i_clk(i_clk));
Mul0000000001  u_000000080C_Mul0000000001(.i_data_1(c_plus_d[171][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[171][2]), .i_clk(i_clk));
Mul0000000001  u_000000080D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[683*12+:12]), .o_data(C[171][2]), .i_clk(i_clk));
Mul0000000001  u_000000080E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[939*12+:12]), .o_data(A[171][3]), .i_clk(i_clk));
Mul0000000001  u_000000080F_Mul0000000001(.i_data_1(c_plus_d[171][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[171][3]), .i_clk(i_clk));
Mul0000000001  u_0000000810_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[939*12+:12]), .o_data(C[171][3]), .i_clk(i_clk));
Mul0000000001  u_0000000811_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[172*12+:12]), .o_data(A[172][0]), .i_clk(i_clk));
Mul0000000001  u_0000000812_Mul0000000001(.i_data_1(c_plus_d[172][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[172][0]), .i_clk(i_clk));
Mul0000000001  u_0000000813_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[172*12+:12]), .o_data(C[172][0]), .i_clk(i_clk));
Mul0000000001  u_0000000814_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[428*12+:12]), .o_data(A[172][1]), .i_clk(i_clk));
Mul0000000001  u_0000000815_Mul0000000001(.i_data_1(c_plus_d[172][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[172][1]), .i_clk(i_clk));
Mul0000000001  u_0000000816_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[428*12+:12]), .o_data(C[172][1]), .i_clk(i_clk));
Mul0000000001  u_0000000817_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[684*12+:12]), .o_data(A[172][2]), .i_clk(i_clk));
Mul0000000001  u_0000000818_Mul0000000001(.i_data_1(c_plus_d[172][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[172][2]), .i_clk(i_clk));
Mul0000000001  u_0000000819_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[684*12+:12]), .o_data(C[172][2]), .i_clk(i_clk));
Mul0000000001  u_000000081A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[940*12+:12]), .o_data(A[172][3]), .i_clk(i_clk));
Mul0000000001  u_000000081B_Mul0000000001(.i_data_1(c_plus_d[172][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[172][3]), .i_clk(i_clk));
Mul0000000001  u_000000081C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[940*12+:12]), .o_data(C[172][3]), .i_clk(i_clk));
Mul0000000001  u_000000081D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[173*12+:12]), .o_data(A[173][0]), .i_clk(i_clk));
Mul0000000001  u_000000081E_Mul0000000001(.i_data_1(c_plus_d[173][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[173][0]), .i_clk(i_clk));
Mul0000000001  u_000000081F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[173*12+:12]), .o_data(C[173][0]), .i_clk(i_clk));
Mul0000000001  u_0000000820_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[429*12+:12]), .o_data(A[173][1]), .i_clk(i_clk));
Mul0000000001  u_0000000821_Mul0000000001(.i_data_1(c_plus_d[173][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[173][1]), .i_clk(i_clk));
Mul0000000001  u_0000000822_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[429*12+:12]), .o_data(C[173][1]), .i_clk(i_clk));
Mul0000000001  u_0000000823_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[685*12+:12]), .o_data(A[173][2]), .i_clk(i_clk));
Mul0000000001  u_0000000824_Mul0000000001(.i_data_1(c_plus_d[173][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[173][2]), .i_clk(i_clk));
Mul0000000001  u_0000000825_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[685*12+:12]), .o_data(C[173][2]), .i_clk(i_clk));
Mul0000000001  u_0000000826_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[941*12+:12]), .o_data(A[173][3]), .i_clk(i_clk));
Mul0000000001  u_0000000827_Mul0000000001(.i_data_1(c_plus_d[173][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[173][3]), .i_clk(i_clk));
Mul0000000001  u_0000000828_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[941*12+:12]), .o_data(C[173][3]), .i_clk(i_clk));
Mul0000000001  u_0000000829_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[174*12+:12]), .o_data(A[174][0]), .i_clk(i_clk));
Mul0000000001  u_000000082A_Mul0000000001(.i_data_1(c_plus_d[174][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[174][0]), .i_clk(i_clk));
Mul0000000001  u_000000082B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[174*12+:12]), .o_data(C[174][0]), .i_clk(i_clk));
Mul0000000001  u_000000082C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[430*12+:12]), .o_data(A[174][1]), .i_clk(i_clk));
Mul0000000001  u_000000082D_Mul0000000001(.i_data_1(c_plus_d[174][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[174][1]), .i_clk(i_clk));
Mul0000000001  u_000000082E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[430*12+:12]), .o_data(C[174][1]), .i_clk(i_clk));
Mul0000000001  u_000000082F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[686*12+:12]), .o_data(A[174][2]), .i_clk(i_clk));
Mul0000000001  u_0000000830_Mul0000000001(.i_data_1(c_plus_d[174][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[174][2]), .i_clk(i_clk));
Mul0000000001  u_0000000831_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[686*12+:12]), .o_data(C[174][2]), .i_clk(i_clk));
Mul0000000001  u_0000000832_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[942*12+:12]), .o_data(A[174][3]), .i_clk(i_clk));
Mul0000000001  u_0000000833_Mul0000000001(.i_data_1(c_plus_d[174][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[174][3]), .i_clk(i_clk));
Mul0000000001  u_0000000834_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[942*12+:12]), .o_data(C[174][3]), .i_clk(i_clk));
Mul0000000001  u_0000000835_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[175*12+:12]), .o_data(A[175][0]), .i_clk(i_clk));
Mul0000000001  u_0000000836_Mul0000000001(.i_data_1(c_plus_d[175][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[175][0]), .i_clk(i_clk));
Mul0000000001  u_0000000837_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[175*12+:12]), .o_data(C[175][0]), .i_clk(i_clk));
Mul0000000001  u_0000000838_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[431*12+:12]), .o_data(A[175][1]), .i_clk(i_clk));
Mul0000000001  u_0000000839_Mul0000000001(.i_data_1(c_plus_d[175][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[175][1]), .i_clk(i_clk));
Mul0000000001  u_000000083A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[431*12+:12]), .o_data(C[175][1]), .i_clk(i_clk));
Mul0000000001  u_000000083B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[687*12+:12]), .o_data(A[175][2]), .i_clk(i_clk));
Mul0000000001  u_000000083C_Mul0000000001(.i_data_1(c_plus_d[175][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[175][2]), .i_clk(i_clk));
Mul0000000001  u_000000083D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[687*12+:12]), .o_data(C[175][2]), .i_clk(i_clk));
Mul0000000001  u_000000083E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[943*12+:12]), .o_data(A[175][3]), .i_clk(i_clk));
Mul0000000001  u_000000083F_Mul0000000001(.i_data_1(c_plus_d[175][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[175][3]), .i_clk(i_clk));
Mul0000000001  u_0000000840_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[943*12+:12]), .o_data(C[175][3]), .i_clk(i_clk));
Mul0000000001  u_0000000841_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[176*12+:12]), .o_data(A[176][0]), .i_clk(i_clk));
Mul0000000001  u_0000000842_Mul0000000001(.i_data_1(c_plus_d[176][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[176][0]), .i_clk(i_clk));
Mul0000000001  u_0000000843_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[176*12+:12]), .o_data(C[176][0]), .i_clk(i_clk));
Mul0000000001  u_0000000844_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[432*12+:12]), .o_data(A[176][1]), .i_clk(i_clk));
Mul0000000001  u_0000000845_Mul0000000001(.i_data_1(c_plus_d[176][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[176][1]), .i_clk(i_clk));
Mul0000000001  u_0000000846_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[432*12+:12]), .o_data(C[176][1]), .i_clk(i_clk));
Mul0000000001  u_0000000847_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[688*12+:12]), .o_data(A[176][2]), .i_clk(i_clk));
Mul0000000001  u_0000000848_Mul0000000001(.i_data_1(c_plus_d[176][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[176][2]), .i_clk(i_clk));
Mul0000000001  u_0000000849_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[688*12+:12]), .o_data(C[176][2]), .i_clk(i_clk));
Mul0000000001  u_000000084A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[944*12+:12]), .o_data(A[176][3]), .i_clk(i_clk));
Mul0000000001  u_000000084B_Mul0000000001(.i_data_1(c_plus_d[176][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[176][3]), .i_clk(i_clk));
Mul0000000001  u_000000084C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[944*12+:12]), .o_data(C[176][3]), .i_clk(i_clk));
Mul0000000001  u_000000084D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[177*12+:12]), .o_data(A[177][0]), .i_clk(i_clk));
Mul0000000001  u_000000084E_Mul0000000001(.i_data_1(c_plus_d[177][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[177][0]), .i_clk(i_clk));
Mul0000000001  u_000000084F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[177*12+:12]), .o_data(C[177][0]), .i_clk(i_clk));
Mul0000000001  u_0000000850_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[433*12+:12]), .o_data(A[177][1]), .i_clk(i_clk));
Mul0000000001  u_0000000851_Mul0000000001(.i_data_1(c_plus_d[177][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[177][1]), .i_clk(i_clk));
Mul0000000001  u_0000000852_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[433*12+:12]), .o_data(C[177][1]), .i_clk(i_clk));
Mul0000000001  u_0000000853_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[689*12+:12]), .o_data(A[177][2]), .i_clk(i_clk));
Mul0000000001  u_0000000854_Mul0000000001(.i_data_1(c_plus_d[177][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[177][2]), .i_clk(i_clk));
Mul0000000001  u_0000000855_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[689*12+:12]), .o_data(C[177][2]), .i_clk(i_clk));
Mul0000000001  u_0000000856_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[945*12+:12]), .o_data(A[177][3]), .i_clk(i_clk));
Mul0000000001  u_0000000857_Mul0000000001(.i_data_1(c_plus_d[177][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[177][3]), .i_clk(i_clk));
Mul0000000001  u_0000000858_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[945*12+:12]), .o_data(C[177][3]), .i_clk(i_clk));
Mul0000000001  u_0000000859_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[178*12+:12]), .o_data(A[178][0]), .i_clk(i_clk));
Mul0000000001  u_000000085A_Mul0000000001(.i_data_1(c_plus_d[178][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[178][0]), .i_clk(i_clk));
Mul0000000001  u_000000085B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[178*12+:12]), .o_data(C[178][0]), .i_clk(i_clk));
Mul0000000001  u_000000085C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[434*12+:12]), .o_data(A[178][1]), .i_clk(i_clk));
Mul0000000001  u_000000085D_Mul0000000001(.i_data_1(c_plus_d[178][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[178][1]), .i_clk(i_clk));
Mul0000000001  u_000000085E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[434*12+:12]), .o_data(C[178][1]), .i_clk(i_clk));
Mul0000000001  u_000000085F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[690*12+:12]), .o_data(A[178][2]), .i_clk(i_clk));
Mul0000000001  u_0000000860_Mul0000000001(.i_data_1(c_plus_d[178][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[178][2]), .i_clk(i_clk));
Mul0000000001  u_0000000861_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[690*12+:12]), .o_data(C[178][2]), .i_clk(i_clk));
Mul0000000001  u_0000000862_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[946*12+:12]), .o_data(A[178][3]), .i_clk(i_clk));
Mul0000000001  u_0000000863_Mul0000000001(.i_data_1(c_plus_d[178][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[178][3]), .i_clk(i_clk));
Mul0000000001  u_0000000864_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[946*12+:12]), .o_data(C[178][3]), .i_clk(i_clk));
Mul0000000001  u_0000000865_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[179*12+:12]), .o_data(A[179][0]), .i_clk(i_clk));
Mul0000000001  u_0000000866_Mul0000000001(.i_data_1(c_plus_d[179][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[179][0]), .i_clk(i_clk));
Mul0000000001  u_0000000867_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[179*12+:12]), .o_data(C[179][0]), .i_clk(i_clk));
Mul0000000001  u_0000000868_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[435*12+:12]), .o_data(A[179][1]), .i_clk(i_clk));
Mul0000000001  u_0000000869_Mul0000000001(.i_data_1(c_plus_d[179][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[179][1]), .i_clk(i_clk));
Mul0000000001  u_000000086A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[435*12+:12]), .o_data(C[179][1]), .i_clk(i_clk));
Mul0000000001  u_000000086B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[691*12+:12]), .o_data(A[179][2]), .i_clk(i_clk));
Mul0000000001  u_000000086C_Mul0000000001(.i_data_1(c_plus_d[179][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[179][2]), .i_clk(i_clk));
Mul0000000001  u_000000086D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[691*12+:12]), .o_data(C[179][2]), .i_clk(i_clk));
Mul0000000001  u_000000086E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[947*12+:12]), .o_data(A[179][3]), .i_clk(i_clk));
Mul0000000001  u_000000086F_Mul0000000001(.i_data_1(c_plus_d[179][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[179][3]), .i_clk(i_clk));
Mul0000000001  u_0000000870_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[947*12+:12]), .o_data(C[179][3]), .i_clk(i_clk));
Mul0000000001  u_0000000871_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[180*12+:12]), .o_data(A[180][0]), .i_clk(i_clk));
Mul0000000001  u_0000000872_Mul0000000001(.i_data_1(c_plus_d[180][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[180][0]), .i_clk(i_clk));
Mul0000000001  u_0000000873_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[180*12+:12]), .o_data(C[180][0]), .i_clk(i_clk));
Mul0000000001  u_0000000874_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[436*12+:12]), .o_data(A[180][1]), .i_clk(i_clk));
Mul0000000001  u_0000000875_Mul0000000001(.i_data_1(c_plus_d[180][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[180][1]), .i_clk(i_clk));
Mul0000000001  u_0000000876_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[436*12+:12]), .o_data(C[180][1]), .i_clk(i_clk));
Mul0000000001  u_0000000877_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[692*12+:12]), .o_data(A[180][2]), .i_clk(i_clk));
Mul0000000001  u_0000000878_Mul0000000001(.i_data_1(c_plus_d[180][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[180][2]), .i_clk(i_clk));
Mul0000000001  u_0000000879_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[692*12+:12]), .o_data(C[180][2]), .i_clk(i_clk));
Mul0000000001  u_000000087A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[948*12+:12]), .o_data(A[180][3]), .i_clk(i_clk));
Mul0000000001  u_000000087B_Mul0000000001(.i_data_1(c_plus_d[180][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[180][3]), .i_clk(i_clk));
Mul0000000001  u_000000087C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[948*12+:12]), .o_data(C[180][3]), .i_clk(i_clk));
Mul0000000001  u_000000087D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[181*12+:12]), .o_data(A[181][0]), .i_clk(i_clk));
Mul0000000001  u_000000087E_Mul0000000001(.i_data_1(c_plus_d[181][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[181][0]), .i_clk(i_clk));
Mul0000000001  u_000000087F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[181*12+:12]), .o_data(C[181][0]), .i_clk(i_clk));
Mul0000000001  u_0000000880_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[437*12+:12]), .o_data(A[181][1]), .i_clk(i_clk));
Mul0000000001  u_0000000881_Mul0000000001(.i_data_1(c_plus_d[181][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[181][1]), .i_clk(i_clk));
Mul0000000001  u_0000000882_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[437*12+:12]), .o_data(C[181][1]), .i_clk(i_clk));
Mul0000000001  u_0000000883_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[693*12+:12]), .o_data(A[181][2]), .i_clk(i_clk));
Mul0000000001  u_0000000884_Mul0000000001(.i_data_1(c_plus_d[181][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[181][2]), .i_clk(i_clk));
Mul0000000001  u_0000000885_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[693*12+:12]), .o_data(C[181][2]), .i_clk(i_clk));
Mul0000000001  u_0000000886_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[949*12+:12]), .o_data(A[181][3]), .i_clk(i_clk));
Mul0000000001  u_0000000887_Mul0000000001(.i_data_1(c_plus_d[181][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[181][3]), .i_clk(i_clk));
Mul0000000001  u_0000000888_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[949*12+:12]), .o_data(C[181][3]), .i_clk(i_clk));
Mul0000000001  u_0000000889_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[182*12+:12]), .o_data(A[182][0]), .i_clk(i_clk));
Mul0000000001  u_000000088A_Mul0000000001(.i_data_1(c_plus_d[182][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[182][0]), .i_clk(i_clk));
Mul0000000001  u_000000088B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[182*12+:12]), .o_data(C[182][0]), .i_clk(i_clk));
Mul0000000001  u_000000088C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[438*12+:12]), .o_data(A[182][1]), .i_clk(i_clk));
Mul0000000001  u_000000088D_Mul0000000001(.i_data_1(c_plus_d[182][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[182][1]), .i_clk(i_clk));
Mul0000000001  u_000000088E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[438*12+:12]), .o_data(C[182][1]), .i_clk(i_clk));
Mul0000000001  u_000000088F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[694*12+:12]), .o_data(A[182][2]), .i_clk(i_clk));
Mul0000000001  u_0000000890_Mul0000000001(.i_data_1(c_plus_d[182][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[182][2]), .i_clk(i_clk));
Mul0000000001  u_0000000891_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[694*12+:12]), .o_data(C[182][2]), .i_clk(i_clk));
Mul0000000001  u_0000000892_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[950*12+:12]), .o_data(A[182][3]), .i_clk(i_clk));
Mul0000000001  u_0000000893_Mul0000000001(.i_data_1(c_plus_d[182][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[182][3]), .i_clk(i_clk));
Mul0000000001  u_0000000894_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[950*12+:12]), .o_data(C[182][3]), .i_clk(i_clk));
Mul0000000001  u_0000000895_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[183*12+:12]), .o_data(A[183][0]), .i_clk(i_clk));
Mul0000000001  u_0000000896_Mul0000000001(.i_data_1(c_plus_d[183][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[183][0]), .i_clk(i_clk));
Mul0000000001  u_0000000897_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[183*12+:12]), .o_data(C[183][0]), .i_clk(i_clk));
Mul0000000001  u_0000000898_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[439*12+:12]), .o_data(A[183][1]), .i_clk(i_clk));
Mul0000000001  u_0000000899_Mul0000000001(.i_data_1(c_plus_d[183][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[183][1]), .i_clk(i_clk));
Mul0000000001  u_000000089A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[439*12+:12]), .o_data(C[183][1]), .i_clk(i_clk));
Mul0000000001  u_000000089B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[695*12+:12]), .o_data(A[183][2]), .i_clk(i_clk));
Mul0000000001  u_000000089C_Mul0000000001(.i_data_1(c_plus_d[183][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[183][2]), .i_clk(i_clk));
Mul0000000001  u_000000089D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[695*12+:12]), .o_data(C[183][2]), .i_clk(i_clk));
Mul0000000001  u_000000089E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[951*12+:12]), .o_data(A[183][3]), .i_clk(i_clk));
Mul0000000001  u_000000089F_Mul0000000001(.i_data_1(c_plus_d[183][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[183][3]), .i_clk(i_clk));
Mul0000000001  u_00000008A0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[951*12+:12]), .o_data(C[183][3]), .i_clk(i_clk));
Mul0000000001  u_00000008A1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[184*12+:12]), .o_data(A[184][0]), .i_clk(i_clk));
Mul0000000001  u_00000008A2_Mul0000000001(.i_data_1(c_plus_d[184][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[184][0]), .i_clk(i_clk));
Mul0000000001  u_00000008A3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[184*12+:12]), .o_data(C[184][0]), .i_clk(i_clk));
Mul0000000001  u_00000008A4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[440*12+:12]), .o_data(A[184][1]), .i_clk(i_clk));
Mul0000000001  u_00000008A5_Mul0000000001(.i_data_1(c_plus_d[184][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[184][1]), .i_clk(i_clk));
Mul0000000001  u_00000008A6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[440*12+:12]), .o_data(C[184][1]), .i_clk(i_clk));
Mul0000000001  u_00000008A7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[696*12+:12]), .o_data(A[184][2]), .i_clk(i_clk));
Mul0000000001  u_00000008A8_Mul0000000001(.i_data_1(c_plus_d[184][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[184][2]), .i_clk(i_clk));
Mul0000000001  u_00000008A9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[696*12+:12]), .o_data(C[184][2]), .i_clk(i_clk));
Mul0000000001  u_00000008AA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[952*12+:12]), .o_data(A[184][3]), .i_clk(i_clk));
Mul0000000001  u_00000008AB_Mul0000000001(.i_data_1(c_plus_d[184][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[184][3]), .i_clk(i_clk));
Mul0000000001  u_00000008AC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[952*12+:12]), .o_data(C[184][3]), .i_clk(i_clk));
Mul0000000001  u_00000008AD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[185*12+:12]), .o_data(A[185][0]), .i_clk(i_clk));
Mul0000000001  u_00000008AE_Mul0000000001(.i_data_1(c_plus_d[185][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[185][0]), .i_clk(i_clk));
Mul0000000001  u_00000008AF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[185*12+:12]), .o_data(C[185][0]), .i_clk(i_clk));
Mul0000000001  u_00000008B0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[441*12+:12]), .o_data(A[185][1]), .i_clk(i_clk));
Mul0000000001  u_00000008B1_Mul0000000001(.i_data_1(c_plus_d[185][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[185][1]), .i_clk(i_clk));
Mul0000000001  u_00000008B2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[441*12+:12]), .o_data(C[185][1]), .i_clk(i_clk));
Mul0000000001  u_00000008B3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[697*12+:12]), .o_data(A[185][2]), .i_clk(i_clk));
Mul0000000001  u_00000008B4_Mul0000000001(.i_data_1(c_plus_d[185][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[185][2]), .i_clk(i_clk));
Mul0000000001  u_00000008B5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[697*12+:12]), .o_data(C[185][2]), .i_clk(i_clk));
Mul0000000001  u_00000008B6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[953*12+:12]), .o_data(A[185][3]), .i_clk(i_clk));
Mul0000000001  u_00000008B7_Mul0000000001(.i_data_1(c_plus_d[185][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[185][3]), .i_clk(i_clk));
Mul0000000001  u_00000008B8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[953*12+:12]), .o_data(C[185][3]), .i_clk(i_clk));
Mul0000000001  u_00000008B9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[186*12+:12]), .o_data(A[186][0]), .i_clk(i_clk));
Mul0000000001  u_00000008BA_Mul0000000001(.i_data_1(c_plus_d[186][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[186][0]), .i_clk(i_clk));
Mul0000000001  u_00000008BB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[186*12+:12]), .o_data(C[186][0]), .i_clk(i_clk));
Mul0000000001  u_00000008BC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[442*12+:12]), .o_data(A[186][1]), .i_clk(i_clk));
Mul0000000001  u_00000008BD_Mul0000000001(.i_data_1(c_plus_d[186][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[186][1]), .i_clk(i_clk));
Mul0000000001  u_00000008BE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[442*12+:12]), .o_data(C[186][1]), .i_clk(i_clk));
Mul0000000001  u_00000008BF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[698*12+:12]), .o_data(A[186][2]), .i_clk(i_clk));
Mul0000000001  u_00000008C0_Mul0000000001(.i_data_1(c_plus_d[186][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[186][2]), .i_clk(i_clk));
Mul0000000001  u_00000008C1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[698*12+:12]), .o_data(C[186][2]), .i_clk(i_clk));
Mul0000000001  u_00000008C2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[954*12+:12]), .o_data(A[186][3]), .i_clk(i_clk));
Mul0000000001  u_00000008C3_Mul0000000001(.i_data_1(c_plus_d[186][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[186][3]), .i_clk(i_clk));
Mul0000000001  u_00000008C4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[954*12+:12]), .o_data(C[186][3]), .i_clk(i_clk));
Mul0000000001  u_00000008C5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[187*12+:12]), .o_data(A[187][0]), .i_clk(i_clk));
Mul0000000001  u_00000008C6_Mul0000000001(.i_data_1(c_plus_d[187][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[187][0]), .i_clk(i_clk));
Mul0000000001  u_00000008C7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[187*12+:12]), .o_data(C[187][0]), .i_clk(i_clk));
Mul0000000001  u_00000008C8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[443*12+:12]), .o_data(A[187][1]), .i_clk(i_clk));
Mul0000000001  u_00000008C9_Mul0000000001(.i_data_1(c_plus_d[187][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[187][1]), .i_clk(i_clk));
Mul0000000001  u_00000008CA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[443*12+:12]), .o_data(C[187][1]), .i_clk(i_clk));
Mul0000000001  u_00000008CB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[699*12+:12]), .o_data(A[187][2]), .i_clk(i_clk));
Mul0000000001  u_00000008CC_Mul0000000001(.i_data_1(c_plus_d[187][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[187][2]), .i_clk(i_clk));
Mul0000000001  u_00000008CD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[699*12+:12]), .o_data(C[187][2]), .i_clk(i_clk));
Mul0000000001  u_00000008CE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[955*12+:12]), .o_data(A[187][3]), .i_clk(i_clk));
Mul0000000001  u_00000008CF_Mul0000000001(.i_data_1(c_plus_d[187][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[187][3]), .i_clk(i_clk));
Mul0000000001  u_00000008D0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[955*12+:12]), .o_data(C[187][3]), .i_clk(i_clk));
Mul0000000001  u_00000008D1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[188*12+:12]), .o_data(A[188][0]), .i_clk(i_clk));
Mul0000000001  u_00000008D2_Mul0000000001(.i_data_1(c_plus_d[188][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[188][0]), .i_clk(i_clk));
Mul0000000001  u_00000008D3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[188*12+:12]), .o_data(C[188][0]), .i_clk(i_clk));
Mul0000000001  u_00000008D4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[444*12+:12]), .o_data(A[188][1]), .i_clk(i_clk));
Mul0000000001  u_00000008D5_Mul0000000001(.i_data_1(c_plus_d[188][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[188][1]), .i_clk(i_clk));
Mul0000000001  u_00000008D6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[444*12+:12]), .o_data(C[188][1]), .i_clk(i_clk));
Mul0000000001  u_00000008D7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[700*12+:12]), .o_data(A[188][2]), .i_clk(i_clk));
Mul0000000001  u_00000008D8_Mul0000000001(.i_data_1(c_plus_d[188][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[188][2]), .i_clk(i_clk));
Mul0000000001  u_00000008D9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[700*12+:12]), .o_data(C[188][2]), .i_clk(i_clk));
Mul0000000001  u_00000008DA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[956*12+:12]), .o_data(A[188][3]), .i_clk(i_clk));
Mul0000000001  u_00000008DB_Mul0000000001(.i_data_1(c_plus_d[188][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[188][3]), .i_clk(i_clk));
Mul0000000001  u_00000008DC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[956*12+:12]), .o_data(C[188][3]), .i_clk(i_clk));
Mul0000000001  u_00000008DD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[189*12+:12]), .o_data(A[189][0]), .i_clk(i_clk));
Mul0000000001  u_00000008DE_Mul0000000001(.i_data_1(c_plus_d[189][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[189][0]), .i_clk(i_clk));
Mul0000000001  u_00000008DF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[189*12+:12]), .o_data(C[189][0]), .i_clk(i_clk));
Mul0000000001  u_00000008E0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[445*12+:12]), .o_data(A[189][1]), .i_clk(i_clk));
Mul0000000001  u_00000008E1_Mul0000000001(.i_data_1(c_plus_d[189][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[189][1]), .i_clk(i_clk));
Mul0000000001  u_00000008E2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[445*12+:12]), .o_data(C[189][1]), .i_clk(i_clk));
Mul0000000001  u_00000008E3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[701*12+:12]), .o_data(A[189][2]), .i_clk(i_clk));
Mul0000000001  u_00000008E4_Mul0000000001(.i_data_1(c_plus_d[189][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[189][2]), .i_clk(i_clk));
Mul0000000001  u_00000008E5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[701*12+:12]), .o_data(C[189][2]), .i_clk(i_clk));
Mul0000000001  u_00000008E6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[957*12+:12]), .o_data(A[189][3]), .i_clk(i_clk));
Mul0000000001  u_00000008E7_Mul0000000001(.i_data_1(c_plus_d[189][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[189][3]), .i_clk(i_clk));
Mul0000000001  u_00000008E8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[957*12+:12]), .o_data(C[189][3]), .i_clk(i_clk));
Mul0000000001  u_00000008E9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[190*12+:12]), .o_data(A[190][0]), .i_clk(i_clk));
Mul0000000001  u_00000008EA_Mul0000000001(.i_data_1(c_plus_d[190][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[190][0]), .i_clk(i_clk));
Mul0000000001  u_00000008EB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[190*12+:12]), .o_data(C[190][0]), .i_clk(i_clk));
Mul0000000001  u_00000008EC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[446*12+:12]), .o_data(A[190][1]), .i_clk(i_clk));
Mul0000000001  u_00000008ED_Mul0000000001(.i_data_1(c_plus_d[190][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[190][1]), .i_clk(i_clk));
Mul0000000001  u_00000008EE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[446*12+:12]), .o_data(C[190][1]), .i_clk(i_clk));
Mul0000000001  u_00000008EF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[702*12+:12]), .o_data(A[190][2]), .i_clk(i_clk));
Mul0000000001  u_00000008F0_Mul0000000001(.i_data_1(c_plus_d[190][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[190][2]), .i_clk(i_clk));
Mul0000000001  u_00000008F1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[702*12+:12]), .o_data(C[190][2]), .i_clk(i_clk));
Mul0000000001  u_00000008F2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[958*12+:12]), .o_data(A[190][3]), .i_clk(i_clk));
Mul0000000001  u_00000008F3_Mul0000000001(.i_data_1(c_plus_d[190][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[190][3]), .i_clk(i_clk));
Mul0000000001  u_00000008F4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[958*12+:12]), .o_data(C[190][3]), .i_clk(i_clk));
Mul0000000001  u_00000008F5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[191*12+:12]), .o_data(A[191][0]), .i_clk(i_clk));
Mul0000000001  u_00000008F6_Mul0000000001(.i_data_1(c_plus_d[191][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[191][0]), .i_clk(i_clk));
Mul0000000001  u_00000008F7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[191*12+:12]), .o_data(C[191][0]), .i_clk(i_clk));
Mul0000000001  u_00000008F8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[447*12+:12]), .o_data(A[191][1]), .i_clk(i_clk));
Mul0000000001  u_00000008F9_Mul0000000001(.i_data_1(c_plus_d[191][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[191][1]), .i_clk(i_clk));
Mul0000000001  u_00000008FA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[447*12+:12]), .o_data(C[191][1]), .i_clk(i_clk));
Mul0000000001  u_00000008FB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[703*12+:12]), .o_data(A[191][2]), .i_clk(i_clk));
Mul0000000001  u_00000008FC_Mul0000000001(.i_data_1(c_plus_d[191][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[191][2]), .i_clk(i_clk));
Mul0000000001  u_00000008FD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[703*12+:12]), .o_data(C[191][2]), .i_clk(i_clk));
Mul0000000001  u_00000008FE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[959*12+:12]), .o_data(A[191][3]), .i_clk(i_clk));
Mul0000000001  u_00000008FF_Mul0000000001(.i_data_1(c_plus_d[191][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[191][3]), .i_clk(i_clk));
Mul0000000001  u_0000000900_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[959*12+:12]), .o_data(C[191][3]), .i_clk(i_clk));
Mul0000000001  u_0000000901_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[192*12+:12]), .o_data(A[192][0]), .i_clk(i_clk));
Mul0000000001  u_0000000902_Mul0000000001(.i_data_1(c_plus_d[192][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[192][0]), .i_clk(i_clk));
Mul0000000001  u_0000000903_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[192*12+:12]), .o_data(C[192][0]), .i_clk(i_clk));
Mul0000000001  u_0000000904_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[448*12+:12]), .o_data(A[192][1]), .i_clk(i_clk));
Mul0000000001  u_0000000905_Mul0000000001(.i_data_1(c_plus_d[192][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[192][1]), .i_clk(i_clk));
Mul0000000001  u_0000000906_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[448*12+:12]), .o_data(C[192][1]), .i_clk(i_clk));
Mul0000000001  u_0000000907_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[704*12+:12]), .o_data(A[192][2]), .i_clk(i_clk));
Mul0000000001  u_0000000908_Mul0000000001(.i_data_1(c_plus_d[192][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[192][2]), .i_clk(i_clk));
Mul0000000001  u_0000000909_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[704*12+:12]), .o_data(C[192][2]), .i_clk(i_clk));
Mul0000000001  u_000000090A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[960*12+:12]), .o_data(A[192][3]), .i_clk(i_clk));
Mul0000000001  u_000000090B_Mul0000000001(.i_data_1(c_plus_d[192][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[192][3]), .i_clk(i_clk));
Mul0000000001  u_000000090C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[960*12+:12]), .o_data(C[192][3]), .i_clk(i_clk));
Mul0000000001  u_000000090D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[193*12+:12]), .o_data(A[193][0]), .i_clk(i_clk));
Mul0000000001  u_000000090E_Mul0000000001(.i_data_1(c_plus_d[193][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[193][0]), .i_clk(i_clk));
Mul0000000001  u_000000090F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[193*12+:12]), .o_data(C[193][0]), .i_clk(i_clk));
Mul0000000001  u_0000000910_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[449*12+:12]), .o_data(A[193][1]), .i_clk(i_clk));
Mul0000000001  u_0000000911_Mul0000000001(.i_data_1(c_plus_d[193][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[193][1]), .i_clk(i_clk));
Mul0000000001  u_0000000912_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[449*12+:12]), .o_data(C[193][1]), .i_clk(i_clk));
Mul0000000001  u_0000000913_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[705*12+:12]), .o_data(A[193][2]), .i_clk(i_clk));
Mul0000000001  u_0000000914_Mul0000000001(.i_data_1(c_plus_d[193][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[193][2]), .i_clk(i_clk));
Mul0000000001  u_0000000915_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[705*12+:12]), .o_data(C[193][2]), .i_clk(i_clk));
Mul0000000001  u_0000000916_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[961*12+:12]), .o_data(A[193][3]), .i_clk(i_clk));
Mul0000000001  u_0000000917_Mul0000000001(.i_data_1(c_plus_d[193][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[193][3]), .i_clk(i_clk));
Mul0000000001  u_0000000918_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[961*12+:12]), .o_data(C[193][3]), .i_clk(i_clk));
Mul0000000001  u_0000000919_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[194*12+:12]), .o_data(A[194][0]), .i_clk(i_clk));
Mul0000000001  u_000000091A_Mul0000000001(.i_data_1(c_plus_d[194][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[194][0]), .i_clk(i_clk));
Mul0000000001  u_000000091B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[194*12+:12]), .o_data(C[194][0]), .i_clk(i_clk));
Mul0000000001  u_000000091C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[450*12+:12]), .o_data(A[194][1]), .i_clk(i_clk));
Mul0000000001  u_000000091D_Mul0000000001(.i_data_1(c_plus_d[194][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[194][1]), .i_clk(i_clk));
Mul0000000001  u_000000091E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[450*12+:12]), .o_data(C[194][1]), .i_clk(i_clk));
Mul0000000001  u_000000091F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[706*12+:12]), .o_data(A[194][2]), .i_clk(i_clk));
Mul0000000001  u_0000000920_Mul0000000001(.i_data_1(c_plus_d[194][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[194][2]), .i_clk(i_clk));
Mul0000000001  u_0000000921_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[706*12+:12]), .o_data(C[194][2]), .i_clk(i_clk));
Mul0000000001  u_0000000922_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[962*12+:12]), .o_data(A[194][3]), .i_clk(i_clk));
Mul0000000001  u_0000000923_Mul0000000001(.i_data_1(c_plus_d[194][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[194][3]), .i_clk(i_clk));
Mul0000000001  u_0000000924_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[962*12+:12]), .o_data(C[194][3]), .i_clk(i_clk));
Mul0000000001  u_0000000925_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[195*12+:12]), .o_data(A[195][0]), .i_clk(i_clk));
Mul0000000001  u_0000000926_Mul0000000001(.i_data_1(c_plus_d[195][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[195][0]), .i_clk(i_clk));
Mul0000000001  u_0000000927_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[195*12+:12]), .o_data(C[195][0]), .i_clk(i_clk));
Mul0000000001  u_0000000928_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[451*12+:12]), .o_data(A[195][1]), .i_clk(i_clk));
Mul0000000001  u_0000000929_Mul0000000001(.i_data_1(c_plus_d[195][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[195][1]), .i_clk(i_clk));
Mul0000000001  u_000000092A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[451*12+:12]), .o_data(C[195][1]), .i_clk(i_clk));
Mul0000000001  u_000000092B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[707*12+:12]), .o_data(A[195][2]), .i_clk(i_clk));
Mul0000000001  u_000000092C_Mul0000000001(.i_data_1(c_plus_d[195][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[195][2]), .i_clk(i_clk));
Mul0000000001  u_000000092D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[707*12+:12]), .o_data(C[195][2]), .i_clk(i_clk));
Mul0000000001  u_000000092E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[963*12+:12]), .o_data(A[195][3]), .i_clk(i_clk));
Mul0000000001  u_000000092F_Mul0000000001(.i_data_1(c_plus_d[195][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[195][3]), .i_clk(i_clk));
Mul0000000001  u_0000000930_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[963*12+:12]), .o_data(C[195][3]), .i_clk(i_clk));
Mul0000000001  u_0000000931_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[196*12+:12]), .o_data(A[196][0]), .i_clk(i_clk));
Mul0000000001  u_0000000932_Mul0000000001(.i_data_1(c_plus_d[196][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[196][0]), .i_clk(i_clk));
Mul0000000001  u_0000000933_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[196*12+:12]), .o_data(C[196][0]), .i_clk(i_clk));
Mul0000000001  u_0000000934_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[452*12+:12]), .o_data(A[196][1]), .i_clk(i_clk));
Mul0000000001  u_0000000935_Mul0000000001(.i_data_1(c_plus_d[196][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[196][1]), .i_clk(i_clk));
Mul0000000001  u_0000000936_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[452*12+:12]), .o_data(C[196][1]), .i_clk(i_clk));
Mul0000000001  u_0000000937_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[708*12+:12]), .o_data(A[196][2]), .i_clk(i_clk));
Mul0000000001  u_0000000938_Mul0000000001(.i_data_1(c_plus_d[196][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[196][2]), .i_clk(i_clk));
Mul0000000001  u_0000000939_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[708*12+:12]), .o_data(C[196][2]), .i_clk(i_clk));
Mul0000000001  u_000000093A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[964*12+:12]), .o_data(A[196][3]), .i_clk(i_clk));
Mul0000000001  u_000000093B_Mul0000000001(.i_data_1(c_plus_d[196][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[196][3]), .i_clk(i_clk));
Mul0000000001  u_000000093C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[964*12+:12]), .o_data(C[196][3]), .i_clk(i_clk));
Mul0000000001  u_000000093D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[197*12+:12]), .o_data(A[197][0]), .i_clk(i_clk));
Mul0000000001  u_000000093E_Mul0000000001(.i_data_1(c_plus_d[197][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[197][0]), .i_clk(i_clk));
Mul0000000001  u_000000093F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[197*12+:12]), .o_data(C[197][0]), .i_clk(i_clk));
Mul0000000001  u_0000000940_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[453*12+:12]), .o_data(A[197][1]), .i_clk(i_clk));
Mul0000000001  u_0000000941_Mul0000000001(.i_data_1(c_plus_d[197][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[197][1]), .i_clk(i_clk));
Mul0000000001  u_0000000942_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[453*12+:12]), .o_data(C[197][1]), .i_clk(i_clk));
Mul0000000001  u_0000000943_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[709*12+:12]), .o_data(A[197][2]), .i_clk(i_clk));
Mul0000000001  u_0000000944_Mul0000000001(.i_data_1(c_plus_d[197][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[197][2]), .i_clk(i_clk));
Mul0000000001  u_0000000945_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[709*12+:12]), .o_data(C[197][2]), .i_clk(i_clk));
Mul0000000001  u_0000000946_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[965*12+:12]), .o_data(A[197][3]), .i_clk(i_clk));
Mul0000000001  u_0000000947_Mul0000000001(.i_data_1(c_plus_d[197][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[197][3]), .i_clk(i_clk));
Mul0000000001  u_0000000948_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[965*12+:12]), .o_data(C[197][3]), .i_clk(i_clk));
Mul0000000001  u_0000000949_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[198*12+:12]), .o_data(A[198][0]), .i_clk(i_clk));
Mul0000000001  u_000000094A_Mul0000000001(.i_data_1(c_plus_d[198][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[198][0]), .i_clk(i_clk));
Mul0000000001  u_000000094B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[198*12+:12]), .o_data(C[198][0]), .i_clk(i_clk));
Mul0000000001  u_000000094C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[454*12+:12]), .o_data(A[198][1]), .i_clk(i_clk));
Mul0000000001  u_000000094D_Mul0000000001(.i_data_1(c_plus_d[198][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[198][1]), .i_clk(i_clk));
Mul0000000001  u_000000094E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[454*12+:12]), .o_data(C[198][1]), .i_clk(i_clk));
Mul0000000001  u_000000094F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[710*12+:12]), .o_data(A[198][2]), .i_clk(i_clk));
Mul0000000001  u_0000000950_Mul0000000001(.i_data_1(c_plus_d[198][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[198][2]), .i_clk(i_clk));
Mul0000000001  u_0000000951_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[710*12+:12]), .o_data(C[198][2]), .i_clk(i_clk));
Mul0000000001  u_0000000952_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[966*12+:12]), .o_data(A[198][3]), .i_clk(i_clk));
Mul0000000001  u_0000000953_Mul0000000001(.i_data_1(c_plus_d[198][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[198][3]), .i_clk(i_clk));
Mul0000000001  u_0000000954_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[966*12+:12]), .o_data(C[198][3]), .i_clk(i_clk));
Mul0000000001  u_0000000955_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[199*12+:12]), .o_data(A[199][0]), .i_clk(i_clk));
Mul0000000001  u_0000000956_Mul0000000001(.i_data_1(c_plus_d[199][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[199][0]), .i_clk(i_clk));
Mul0000000001  u_0000000957_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[199*12+:12]), .o_data(C[199][0]), .i_clk(i_clk));
Mul0000000001  u_0000000958_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[455*12+:12]), .o_data(A[199][1]), .i_clk(i_clk));
Mul0000000001  u_0000000959_Mul0000000001(.i_data_1(c_plus_d[199][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[199][1]), .i_clk(i_clk));
Mul0000000001  u_000000095A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[455*12+:12]), .o_data(C[199][1]), .i_clk(i_clk));
Mul0000000001  u_000000095B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[711*12+:12]), .o_data(A[199][2]), .i_clk(i_clk));
Mul0000000001  u_000000095C_Mul0000000001(.i_data_1(c_plus_d[199][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[199][2]), .i_clk(i_clk));
Mul0000000001  u_000000095D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[711*12+:12]), .o_data(C[199][2]), .i_clk(i_clk));
Mul0000000001  u_000000095E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[967*12+:12]), .o_data(A[199][3]), .i_clk(i_clk));
Mul0000000001  u_000000095F_Mul0000000001(.i_data_1(c_plus_d[199][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[199][3]), .i_clk(i_clk));
Mul0000000001  u_0000000960_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[967*12+:12]), .o_data(C[199][3]), .i_clk(i_clk));
Mul0000000001  u_0000000961_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[200*12+:12]), .o_data(A[200][0]), .i_clk(i_clk));
Mul0000000001  u_0000000962_Mul0000000001(.i_data_1(c_plus_d[200][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[200][0]), .i_clk(i_clk));
Mul0000000001  u_0000000963_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[200*12+:12]), .o_data(C[200][0]), .i_clk(i_clk));
Mul0000000001  u_0000000964_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[456*12+:12]), .o_data(A[200][1]), .i_clk(i_clk));
Mul0000000001  u_0000000965_Mul0000000001(.i_data_1(c_plus_d[200][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[200][1]), .i_clk(i_clk));
Mul0000000001  u_0000000966_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[456*12+:12]), .o_data(C[200][1]), .i_clk(i_clk));
Mul0000000001  u_0000000967_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[712*12+:12]), .o_data(A[200][2]), .i_clk(i_clk));
Mul0000000001  u_0000000968_Mul0000000001(.i_data_1(c_plus_d[200][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[200][2]), .i_clk(i_clk));
Mul0000000001  u_0000000969_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[712*12+:12]), .o_data(C[200][2]), .i_clk(i_clk));
Mul0000000001  u_000000096A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[968*12+:12]), .o_data(A[200][3]), .i_clk(i_clk));
Mul0000000001  u_000000096B_Mul0000000001(.i_data_1(c_plus_d[200][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[200][3]), .i_clk(i_clk));
Mul0000000001  u_000000096C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[968*12+:12]), .o_data(C[200][3]), .i_clk(i_clk));
Mul0000000001  u_000000096D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[201*12+:12]), .o_data(A[201][0]), .i_clk(i_clk));
Mul0000000001  u_000000096E_Mul0000000001(.i_data_1(c_plus_d[201][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[201][0]), .i_clk(i_clk));
Mul0000000001  u_000000096F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[201*12+:12]), .o_data(C[201][0]), .i_clk(i_clk));
Mul0000000001  u_0000000970_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[457*12+:12]), .o_data(A[201][1]), .i_clk(i_clk));
Mul0000000001  u_0000000971_Mul0000000001(.i_data_1(c_plus_d[201][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[201][1]), .i_clk(i_clk));
Mul0000000001  u_0000000972_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[457*12+:12]), .o_data(C[201][1]), .i_clk(i_clk));
Mul0000000001  u_0000000973_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[713*12+:12]), .o_data(A[201][2]), .i_clk(i_clk));
Mul0000000001  u_0000000974_Mul0000000001(.i_data_1(c_plus_d[201][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[201][2]), .i_clk(i_clk));
Mul0000000001  u_0000000975_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[713*12+:12]), .o_data(C[201][2]), .i_clk(i_clk));
Mul0000000001  u_0000000976_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[969*12+:12]), .o_data(A[201][3]), .i_clk(i_clk));
Mul0000000001  u_0000000977_Mul0000000001(.i_data_1(c_plus_d[201][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[201][3]), .i_clk(i_clk));
Mul0000000001  u_0000000978_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[969*12+:12]), .o_data(C[201][3]), .i_clk(i_clk));
Mul0000000001  u_0000000979_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[202*12+:12]), .o_data(A[202][0]), .i_clk(i_clk));
Mul0000000001  u_000000097A_Mul0000000001(.i_data_1(c_plus_d[202][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[202][0]), .i_clk(i_clk));
Mul0000000001  u_000000097B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[202*12+:12]), .o_data(C[202][0]), .i_clk(i_clk));
Mul0000000001  u_000000097C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[458*12+:12]), .o_data(A[202][1]), .i_clk(i_clk));
Mul0000000001  u_000000097D_Mul0000000001(.i_data_1(c_plus_d[202][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[202][1]), .i_clk(i_clk));
Mul0000000001  u_000000097E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[458*12+:12]), .o_data(C[202][1]), .i_clk(i_clk));
Mul0000000001  u_000000097F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[714*12+:12]), .o_data(A[202][2]), .i_clk(i_clk));
Mul0000000001  u_0000000980_Mul0000000001(.i_data_1(c_plus_d[202][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[202][2]), .i_clk(i_clk));
Mul0000000001  u_0000000981_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[714*12+:12]), .o_data(C[202][2]), .i_clk(i_clk));
Mul0000000001  u_0000000982_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[970*12+:12]), .o_data(A[202][3]), .i_clk(i_clk));
Mul0000000001  u_0000000983_Mul0000000001(.i_data_1(c_plus_d[202][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[202][3]), .i_clk(i_clk));
Mul0000000001  u_0000000984_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[970*12+:12]), .o_data(C[202][3]), .i_clk(i_clk));
Mul0000000001  u_0000000985_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[203*12+:12]), .o_data(A[203][0]), .i_clk(i_clk));
Mul0000000001  u_0000000986_Mul0000000001(.i_data_1(c_plus_d[203][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[203][0]), .i_clk(i_clk));
Mul0000000001  u_0000000987_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[203*12+:12]), .o_data(C[203][0]), .i_clk(i_clk));
Mul0000000001  u_0000000988_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[459*12+:12]), .o_data(A[203][1]), .i_clk(i_clk));
Mul0000000001  u_0000000989_Mul0000000001(.i_data_1(c_plus_d[203][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[203][1]), .i_clk(i_clk));
Mul0000000001  u_000000098A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[459*12+:12]), .o_data(C[203][1]), .i_clk(i_clk));
Mul0000000001  u_000000098B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[715*12+:12]), .o_data(A[203][2]), .i_clk(i_clk));
Mul0000000001  u_000000098C_Mul0000000001(.i_data_1(c_plus_d[203][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[203][2]), .i_clk(i_clk));
Mul0000000001  u_000000098D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[715*12+:12]), .o_data(C[203][2]), .i_clk(i_clk));
Mul0000000001  u_000000098E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[971*12+:12]), .o_data(A[203][3]), .i_clk(i_clk));
Mul0000000001  u_000000098F_Mul0000000001(.i_data_1(c_plus_d[203][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[203][3]), .i_clk(i_clk));
Mul0000000001  u_0000000990_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[971*12+:12]), .o_data(C[203][3]), .i_clk(i_clk));
Mul0000000001  u_0000000991_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[204*12+:12]), .o_data(A[204][0]), .i_clk(i_clk));
Mul0000000001  u_0000000992_Mul0000000001(.i_data_1(c_plus_d[204][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[204][0]), .i_clk(i_clk));
Mul0000000001  u_0000000993_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[204*12+:12]), .o_data(C[204][0]), .i_clk(i_clk));
Mul0000000001  u_0000000994_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[460*12+:12]), .o_data(A[204][1]), .i_clk(i_clk));
Mul0000000001  u_0000000995_Mul0000000001(.i_data_1(c_plus_d[204][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[204][1]), .i_clk(i_clk));
Mul0000000001  u_0000000996_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[460*12+:12]), .o_data(C[204][1]), .i_clk(i_clk));
Mul0000000001  u_0000000997_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[716*12+:12]), .o_data(A[204][2]), .i_clk(i_clk));
Mul0000000001  u_0000000998_Mul0000000001(.i_data_1(c_plus_d[204][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[204][2]), .i_clk(i_clk));
Mul0000000001  u_0000000999_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[716*12+:12]), .o_data(C[204][2]), .i_clk(i_clk));
Mul0000000001  u_000000099A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[972*12+:12]), .o_data(A[204][3]), .i_clk(i_clk));
Mul0000000001  u_000000099B_Mul0000000001(.i_data_1(c_plus_d[204][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[204][3]), .i_clk(i_clk));
Mul0000000001  u_000000099C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[972*12+:12]), .o_data(C[204][3]), .i_clk(i_clk));
Mul0000000001  u_000000099D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[205*12+:12]), .o_data(A[205][0]), .i_clk(i_clk));
Mul0000000001  u_000000099E_Mul0000000001(.i_data_1(c_plus_d[205][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[205][0]), .i_clk(i_clk));
Mul0000000001  u_000000099F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[205*12+:12]), .o_data(C[205][0]), .i_clk(i_clk));
Mul0000000001  u_00000009A0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[461*12+:12]), .o_data(A[205][1]), .i_clk(i_clk));
Mul0000000001  u_00000009A1_Mul0000000001(.i_data_1(c_plus_d[205][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[205][1]), .i_clk(i_clk));
Mul0000000001  u_00000009A2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[461*12+:12]), .o_data(C[205][1]), .i_clk(i_clk));
Mul0000000001  u_00000009A3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[717*12+:12]), .o_data(A[205][2]), .i_clk(i_clk));
Mul0000000001  u_00000009A4_Mul0000000001(.i_data_1(c_plus_d[205][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[205][2]), .i_clk(i_clk));
Mul0000000001  u_00000009A5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[717*12+:12]), .o_data(C[205][2]), .i_clk(i_clk));
Mul0000000001  u_00000009A6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[973*12+:12]), .o_data(A[205][3]), .i_clk(i_clk));
Mul0000000001  u_00000009A7_Mul0000000001(.i_data_1(c_plus_d[205][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[205][3]), .i_clk(i_clk));
Mul0000000001  u_00000009A8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[973*12+:12]), .o_data(C[205][3]), .i_clk(i_clk));
Mul0000000001  u_00000009A9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[206*12+:12]), .o_data(A[206][0]), .i_clk(i_clk));
Mul0000000001  u_00000009AA_Mul0000000001(.i_data_1(c_plus_d[206][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[206][0]), .i_clk(i_clk));
Mul0000000001  u_00000009AB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[206*12+:12]), .o_data(C[206][0]), .i_clk(i_clk));
Mul0000000001  u_00000009AC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[462*12+:12]), .o_data(A[206][1]), .i_clk(i_clk));
Mul0000000001  u_00000009AD_Mul0000000001(.i_data_1(c_plus_d[206][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[206][1]), .i_clk(i_clk));
Mul0000000001  u_00000009AE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[462*12+:12]), .o_data(C[206][1]), .i_clk(i_clk));
Mul0000000001  u_00000009AF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[718*12+:12]), .o_data(A[206][2]), .i_clk(i_clk));
Mul0000000001  u_00000009B0_Mul0000000001(.i_data_1(c_plus_d[206][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[206][2]), .i_clk(i_clk));
Mul0000000001  u_00000009B1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[718*12+:12]), .o_data(C[206][2]), .i_clk(i_clk));
Mul0000000001  u_00000009B2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[974*12+:12]), .o_data(A[206][3]), .i_clk(i_clk));
Mul0000000001  u_00000009B3_Mul0000000001(.i_data_1(c_plus_d[206][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[206][3]), .i_clk(i_clk));
Mul0000000001  u_00000009B4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[974*12+:12]), .o_data(C[206][3]), .i_clk(i_clk));
Mul0000000001  u_00000009B5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[207*12+:12]), .o_data(A[207][0]), .i_clk(i_clk));
Mul0000000001  u_00000009B6_Mul0000000001(.i_data_1(c_plus_d[207][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[207][0]), .i_clk(i_clk));
Mul0000000001  u_00000009B7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[207*12+:12]), .o_data(C[207][0]), .i_clk(i_clk));
Mul0000000001  u_00000009B8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[463*12+:12]), .o_data(A[207][1]), .i_clk(i_clk));
Mul0000000001  u_00000009B9_Mul0000000001(.i_data_1(c_plus_d[207][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[207][1]), .i_clk(i_clk));
Mul0000000001  u_00000009BA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[463*12+:12]), .o_data(C[207][1]), .i_clk(i_clk));
Mul0000000001  u_00000009BB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[719*12+:12]), .o_data(A[207][2]), .i_clk(i_clk));
Mul0000000001  u_00000009BC_Mul0000000001(.i_data_1(c_plus_d[207][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[207][2]), .i_clk(i_clk));
Mul0000000001  u_00000009BD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[719*12+:12]), .o_data(C[207][2]), .i_clk(i_clk));
Mul0000000001  u_00000009BE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[975*12+:12]), .o_data(A[207][3]), .i_clk(i_clk));
Mul0000000001  u_00000009BF_Mul0000000001(.i_data_1(c_plus_d[207][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[207][3]), .i_clk(i_clk));
Mul0000000001  u_00000009C0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[975*12+:12]), .o_data(C[207][3]), .i_clk(i_clk));
Mul0000000001  u_00000009C1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[208*12+:12]), .o_data(A[208][0]), .i_clk(i_clk));
Mul0000000001  u_00000009C2_Mul0000000001(.i_data_1(c_plus_d[208][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[208][0]), .i_clk(i_clk));
Mul0000000001  u_00000009C3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[208*12+:12]), .o_data(C[208][0]), .i_clk(i_clk));
Mul0000000001  u_00000009C4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[464*12+:12]), .o_data(A[208][1]), .i_clk(i_clk));
Mul0000000001  u_00000009C5_Mul0000000001(.i_data_1(c_plus_d[208][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[208][1]), .i_clk(i_clk));
Mul0000000001  u_00000009C6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[464*12+:12]), .o_data(C[208][1]), .i_clk(i_clk));
Mul0000000001  u_00000009C7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[720*12+:12]), .o_data(A[208][2]), .i_clk(i_clk));
Mul0000000001  u_00000009C8_Mul0000000001(.i_data_1(c_plus_d[208][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[208][2]), .i_clk(i_clk));
Mul0000000001  u_00000009C9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[720*12+:12]), .o_data(C[208][2]), .i_clk(i_clk));
Mul0000000001  u_00000009CA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[976*12+:12]), .o_data(A[208][3]), .i_clk(i_clk));
Mul0000000001  u_00000009CB_Mul0000000001(.i_data_1(c_plus_d[208][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[208][3]), .i_clk(i_clk));
Mul0000000001  u_00000009CC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[976*12+:12]), .o_data(C[208][3]), .i_clk(i_clk));
Mul0000000001  u_00000009CD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[209*12+:12]), .o_data(A[209][0]), .i_clk(i_clk));
Mul0000000001  u_00000009CE_Mul0000000001(.i_data_1(c_plus_d[209][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[209][0]), .i_clk(i_clk));
Mul0000000001  u_00000009CF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[209*12+:12]), .o_data(C[209][0]), .i_clk(i_clk));
Mul0000000001  u_00000009D0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[465*12+:12]), .o_data(A[209][1]), .i_clk(i_clk));
Mul0000000001  u_00000009D1_Mul0000000001(.i_data_1(c_plus_d[209][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[209][1]), .i_clk(i_clk));
Mul0000000001  u_00000009D2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[465*12+:12]), .o_data(C[209][1]), .i_clk(i_clk));
Mul0000000001  u_00000009D3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[721*12+:12]), .o_data(A[209][2]), .i_clk(i_clk));
Mul0000000001  u_00000009D4_Mul0000000001(.i_data_1(c_plus_d[209][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[209][2]), .i_clk(i_clk));
Mul0000000001  u_00000009D5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[721*12+:12]), .o_data(C[209][2]), .i_clk(i_clk));
Mul0000000001  u_00000009D6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[977*12+:12]), .o_data(A[209][3]), .i_clk(i_clk));
Mul0000000001  u_00000009D7_Mul0000000001(.i_data_1(c_plus_d[209][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[209][3]), .i_clk(i_clk));
Mul0000000001  u_00000009D8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[977*12+:12]), .o_data(C[209][3]), .i_clk(i_clk));
Mul0000000001  u_00000009D9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[210*12+:12]), .o_data(A[210][0]), .i_clk(i_clk));
Mul0000000001  u_00000009DA_Mul0000000001(.i_data_1(c_plus_d[210][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[210][0]), .i_clk(i_clk));
Mul0000000001  u_00000009DB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[210*12+:12]), .o_data(C[210][0]), .i_clk(i_clk));
Mul0000000001  u_00000009DC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[466*12+:12]), .o_data(A[210][1]), .i_clk(i_clk));
Mul0000000001  u_00000009DD_Mul0000000001(.i_data_1(c_plus_d[210][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[210][1]), .i_clk(i_clk));
Mul0000000001  u_00000009DE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[466*12+:12]), .o_data(C[210][1]), .i_clk(i_clk));
Mul0000000001  u_00000009DF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[722*12+:12]), .o_data(A[210][2]), .i_clk(i_clk));
Mul0000000001  u_00000009E0_Mul0000000001(.i_data_1(c_plus_d[210][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[210][2]), .i_clk(i_clk));
Mul0000000001  u_00000009E1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[722*12+:12]), .o_data(C[210][2]), .i_clk(i_clk));
Mul0000000001  u_00000009E2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[978*12+:12]), .o_data(A[210][3]), .i_clk(i_clk));
Mul0000000001  u_00000009E3_Mul0000000001(.i_data_1(c_plus_d[210][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[210][3]), .i_clk(i_clk));
Mul0000000001  u_00000009E4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[978*12+:12]), .o_data(C[210][3]), .i_clk(i_clk));
Mul0000000001  u_00000009E5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[211*12+:12]), .o_data(A[211][0]), .i_clk(i_clk));
Mul0000000001  u_00000009E6_Mul0000000001(.i_data_1(c_plus_d[211][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[211][0]), .i_clk(i_clk));
Mul0000000001  u_00000009E7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[211*12+:12]), .o_data(C[211][0]), .i_clk(i_clk));
Mul0000000001  u_00000009E8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[467*12+:12]), .o_data(A[211][1]), .i_clk(i_clk));
Mul0000000001  u_00000009E9_Mul0000000001(.i_data_1(c_plus_d[211][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[211][1]), .i_clk(i_clk));
Mul0000000001  u_00000009EA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[467*12+:12]), .o_data(C[211][1]), .i_clk(i_clk));
Mul0000000001  u_00000009EB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[723*12+:12]), .o_data(A[211][2]), .i_clk(i_clk));
Mul0000000001  u_00000009EC_Mul0000000001(.i_data_1(c_plus_d[211][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[211][2]), .i_clk(i_clk));
Mul0000000001  u_00000009ED_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[723*12+:12]), .o_data(C[211][2]), .i_clk(i_clk));
Mul0000000001  u_00000009EE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[979*12+:12]), .o_data(A[211][3]), .i_clk(i_clk));
Mul0000000001  u_00000009EF_Mul0000000001(.i_data_1(c_plus_d[211][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[211][3]), .i_clk(i_clk));
Mul0000000001  u_00000009F0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[979*12+:12]), .o_data(C[211][3]), .i_clk(i_clk));
Mul0000000001  u_00000009F1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[212*12+:12]), .o_data(A[212][0]), .i_clk(i_clk));
Mul0000000001  u_00000009F2_Mul0000000001(.i_data_1(c_plus_d[212][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[212][0]), .i_clk(i_clk));
Mul0000000001  u_00000009F3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[212*12+:12]), .o_data(C[212][0]), .i_clk(i_clk));
Mul0000000001  u_00000009F4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[468*12+:12]), .o_data(A[212][1]), .i_clk(i_clk));
Mul0000000001  u_00000009F5_Mul0000000001(.i_data_1(c_plus_d[212][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[212][1]), .i_clk(i_clk));
Mul0000000001  u_00000009F6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[468*12+:12]), .o_data(C[212][1]), .i_clk(i_clk));
Mul0000000001  u_00000009F7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[724*12+:12]), .o_data(A[212][2]), .i_clk(i_clk));
Mul0000000001  u_00000009F8_Mul0000000001(.i_data_1(c_plus_d[212][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[212][2]), .i_clk(i_clk));
Mul0000000001  u_00000009F9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[724*12+:12]), .o_data(C[212][2]), .i_clk(i_clk));
Mul0000000001  u_00000009FA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[980*12+:12]), .o_data(A[212][3]), .i_clk(i_clk));
Mul0000000001  u_00000009FB_Mul0000000001(.i_data_1(c_plus_d[212][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[212][3]), .i_clk(i_clk));
Mul0000000001  u_00000009FC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[980*12+:12]), .o_data(C[212][3]), .i_clk(i_clk));
Mul0000000001  u_00000009FD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[213*12+:12]), .o_data(A[213][0]), .i_clk(i_clk));
Mul0000000001  u_00000009FE_Mul0000000001(.i_data_1(c_plus_d[213][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[213][0]), .i_clk(i_clk));
Mul0000000001  u_00000009FF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[213*12+:12]), .o_data(C[213][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A00_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[469*12+:12]), .o_data(A[213][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A01_Mul0000000001(.i_data_1(c_plus_d[213][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[213][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A02_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[469*12+:12]), .o_data(C[213][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A03_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[725*12+:12]), .o_data(A[213][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A04_Mul0000000001(.i_data_1(c_plus_d[213][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[213][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A05_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[725*12+:12]), .o_data(C[213][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A06_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[981*12+:12]), .o_data(A[213][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A07_Mul0000000001(.i_data_1(c_plus_d[213][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[213][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A08_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[981*12+:12]), .o_data(C[213][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A09_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[214*12+:12]), .o_data(A[214][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A0A_Mul0000000001(.i_data_1(c_plus_d[214][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[214][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A0B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[214*12+:12]), .o_data(C[214][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A0C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[470*12+:12]), .o_data(A[214][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A0D_Mul0000000001(.i_data_1(c_plus_d[214][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[214][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A0E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[470*12+:12]), .o_data(C[214][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A0F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[726*12+:12]), .o_data(A[214][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A10_Mul0000000001(.i_data_1(c_plus_d[214][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[214][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A11_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[726*12+:12]), .o_data(C[214][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A12_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[982*12+:12]), .o_data(A[214][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A13_Mul0000000001(.i_data_1(c_plus_d[214][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[214][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A14_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[982*12+:12]), .o_data(C[214][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A15_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[215*12+:12]), .o_data(A[215][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A16_Mul0000000001(.i_data_1(c_plus_d[215][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[215][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A17_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[215*12+:12]), .o_data(C[215][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A18_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[471*12+:12]), .o_data(A[215][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A19_Mul0000000001(.i_data_1(c_plus_d[215][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[215][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A1A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[471*12+:12]), .o_data(C[215][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A1B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[727*12+:12]), .o_data(A[215][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A1C_Mul0000000001(.i_data_1(c_plus_d[215][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[215][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A1D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[727*12+:12]), .o_data(C[215][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A1E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[983*12+:12]), .o_data(A[215][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A1F_Mul0000000001(.i_data_1(c_plus_d[215][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[215][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A20_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[983*12+:12]), .o_data(C[215][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A21_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[216*12+:12]), .o_data(A[216][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A22_Mul0000000001(.i_data_1(c_plus_d[216][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[216][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A23_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[216*12+:12]), .o_data(C[216][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A24_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[472*12+:12]), .o_data(A[216][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A25_Mul0000000001(.i_data_1(c_plus_d[216][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[216][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A26_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[472*12+:12]), .o_data(C[216][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A27_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[728*12+:12]), .o_data(A[216][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A28_Mul0000000001(.i_data_1(c_plus_d[216][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[216][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A29_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[728*12+:12]), .o_data(C[216][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A2A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[984*12+:12]), .o_data(A[216][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A2B_Mul0000000001(.i_data_1(c_plus_d[216][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[216][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A2C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[984*12+:12]), .o_data(C[216][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A2D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[217*12+:12]), .o_data(A[217][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A2E_Mul0000000001(.i_data_1(c_plus_d[217][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[217][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A2F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[217*12+:12]), .o_data(C[217][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A30_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[473*12+:12]), .o_data(A[217][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A31_Mul0000000001(.i_data_1(c_plus_d[217][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[217][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A32_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[473*12+:12]), .o_data(C[217][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A33_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[729*12+:12]), .o_data(A[217][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A34_Mul0000000001(.i_data_1(c_plus_d[217][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[217][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A35_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[729*12+:12]), .o_data(C[217][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A36_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[985*12+:12]), .o_data(A[217][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A37_Mul0000000001(.i_data_1(c_plus_d[217][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[217][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A38_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[985*12+:12]), .o_data(C[217][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A39_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[218*12+:12]), .o_data(A[218][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A3A_Mul0000000001(.i_data_1(c_plus_d[218][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[218][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A3B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[218*12+:12]), .o_data(C[218][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A3C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[474*12+:12]), .o_data(A[218][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A3D_Mul0000000001(.i_data_1(c_plus_d[218][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[218][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A3E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[474*12+:12]), .o_data(C[218][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A3F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[730*12+:12]), .o_data(A[218][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A40_Mul0000000001(.i_data_1(c_plus_d[218][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[218][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A41_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[730*12+:12]), .o_data(C[218][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A42_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[986*12+:12]), .o_data(A[218][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A43_Mul0000000001(.i_data_1(c_plus_d[218][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[218][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A44_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[986*12+:12]), .o_data(C[218][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A45_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[219*12+:12]), .o_data(A[219][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A46_Mul0000000001(.i_data_1(c_plus_d[219][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[219][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A47_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[219*12+:12]), .o_data(C[219][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A48_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[475*12+:12]), .o_data(A[219][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A49_Mul0000000001(.i_data_1(c_plus_d[219][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[219][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A4A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[475*12+:12]), .o_data(C[219][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A4B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[731*12+:12]), .o_data(A[219][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A4C_Mul0000000001(.i_data_1(c_plus_d[219][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[219][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A4D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[731*12+:12]), .o_data(C[219][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A4E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[987*12+:12]), .o_data(A[219][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A4F_Mul0000000001(.i_data_1(c_plus_d[219][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[219][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A50_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[987*12+:12]), .o_data(C[219][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A51_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[220*12+:12]), .o_data(A[220][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A52_Mul0000000001(.i_data_1(c_plus_d[220][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[220][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A53_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[220*12+:12]), .o_data(C[220][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A54_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[476*12+:12]), .o_data(A[220][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A55_Mul0000000001(.i_data_1(c_plus_d[220][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[220][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A56_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[476*12+:12]), .o_data(C[220][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A57_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[732*12+:12]), .o_data(A[220][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A58_Mul0000000001(.i_data_1(c_plus_d[220][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[220][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A59_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[732*12+:12]), .o_data(C[220][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A5A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[988*12+:12]), .o_data(A[220][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A5B_Mul0000000001(.i_data_1(c_plus_d[220][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[220][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A5C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[988*12+:12]), .o_data(C[220][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A5D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[221*12+:12]), .o_data(A[221][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A5E_Mul0000000001(.i_data_1(c_plus_d[221][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[221][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A5F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[221*12+:12]), .o_data(C[221][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A60_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[477*12+:12]), .o_data(A[221][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A61_Mul0000000001(.i_data_1(c_plus_d[221][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[221][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A62_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[477*12+:12]), .o_data(C[221][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A63_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[733*12+:12]), .o_data(A[221][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A64_Mul0000000001(.i_data_1(c_plus_d[221][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[221][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A65_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[733*12+:12]), .o_data(C[221][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A66_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[989*12+:12]), .o_data(A[221][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A67_Mul0000000001(.i_data_1(c_plus_d[221][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[221][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A68_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[989*12+:12]), .o_data(C[221][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A69_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[222*12+:12]), .o_data(A[222][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A6A_Mul0000000001(.i_data_1(c_plus_d[222][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[222][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A6B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[222*12+:12]), .o_data(C[222][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A6C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[478*12+:12]), .o_data(A[222][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A6D_Mul0000000001(.i_data_1(c_plus_d[222][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[222][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A6E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[478*12+:12]), .o_data(C[222][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A6F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[734*12+:12]), .o_data(A[222][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A70_Mul0000000001(.i_data_1(c_plus_d[222][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[222][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A71_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[734*12+:12]), .o_data(C[222][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A72_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[990*12+:12]), .o_data(A[222][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A73_Mul0000000001(.i_data_1(c_plus_d[222][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[222][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A74_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[990*12+:12]), .o_data(C[222][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A75_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[223*12+:12]), .o_data(A[223][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A76_Mul0000000001(.i_data_1(c_plus_d[223][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[223][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A77_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[223*12+:12]), .o_data(C[223][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A78_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[479*12+:12]), .o_data(A[223][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A79_Mul0000000001(.i_data_1(c_plus_d[223][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[223][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A7A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[479*12+:12]), .o_data(C[223][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A7B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[735*12+:12]), .o_data(A[223][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A7C_Mul0000000001(.i_data_1(c_plus_d[223][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[223][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A7D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[735*12+:12]), .o_data(C[223][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A7E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[991*12+:12]), .o_data(A[223][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A7F_Mul0000000001(.i_data_1(c_plus_d[223][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[223][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A80_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[991*12+:12]), .o_data(C[223][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A81_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[224*12+:12]), .o_data(A[224][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A82_Mul0000000001(.i_data_1(c_plus_d[224][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[224][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A83_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[224*12+:12]), .o_data(C[224][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A84_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[480*12+:12]), .o_data(A[224][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A85_Mul0000000001(.i_data_1(c_plus_d[224][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[224][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A86_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[480*12+:12]), .o_data(C[224][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A87_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[736*12+:12]), .o_data(A[224][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A88_Mul0000000001(.i_data_1(c_plus_d[224][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[224][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A89_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[736*12+:12]), .o_data(C[224][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A8A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[992*12+:12]), .o_data(A[224][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A8B_Mul0000000001(.i_data_1(c_plus_d[224][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[224][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A8C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[992*12+:12]), .o_data(C[224][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A8D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[225*12+:12]), .o_data(A[225][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A8E_Mul0000000001(.i_data_1(c_plus_d[225][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[225][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A8F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[225*12+:12]), .o_data(C[225][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A90_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[481*12+:12]), .o_data(A[225][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A91_Mul0000000001(.i_data_1(c_plus_d[225][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[225][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A92_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[481*12+:12]), .o_data(C[225][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A93_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[737*12+:12]), .o_data(A[225][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A94_Mul0000000001(.i_data_1(c_plus_d[225][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[225][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A95_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[737*12+:12]), .o_data(C[225][2]), .i_clk(i_clk));
Mul0000000001  u_0000000A96_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[993*12+:12]), .o_data(A[225][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A97_Mul0000000001(.i_data_1(c_plus_d[225][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[225][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A98_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[993*12+:12]), .o_data(C[225][3]), .i_clk(i_clk));
Mul0000000001  u_0000000A99_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[226*12+:12]), .o_data(A[226][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A9A_Mul0000000001(.i_data_1(c_plus_d[226][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[226][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A9B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[226*12+:12]), .o_data(C[226][0]), .i_clk(i_clk));
Mul0000000001  u_0000000A9C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[482*12+:12]), .o_data(A[226][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A9D_Mul0000000001(.i_data_1(c_plus_d[226][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[226][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A9E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[482*12+:12]), .o_data(C[226][1]), .i_clk(i_clk));
Mul0000000001  u_0000000A9F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[738*12+:12]), .o_data(A[226][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AA0_Mul0000000001(.i_data_1(c_plus_d[226][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[226][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AA1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[738*12+:12]), .o_data(C[226][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AA2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[994*12+:12]), .o_data(A[226][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AA3_Mul0000000001(.i_data_1(c_plus_d[226][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[226][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AA4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[994*12+:12]), .o_data(C[226][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AA5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[227*12+:12]), .o_data(A[227][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AA6_Mul0000000001(.i_data_1(c_plus_d[227][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[227][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AA7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[227*12+:12]), .o_data(C[227][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AA8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[483*12+:12]), .o_data(A[227][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AA9_Mul0000000001(.i_data_1(c_plus_d[227][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[227][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AAA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[483*12+:12]), .o_data(C[227][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AAB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[739*12+:12]), .o_data(A[227][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AAC_Mul0000000001(.i_data_1(c_plus_d[227][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[227][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AAD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[739*12+:12]), .o_data(C[227][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AAE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[995*12+:12]), .o_data(A[227][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AAF_Mul0000000001(.i_data_1(c_plus_d[227][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[227][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AB0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[995*12+:12]), .o_data(C[227][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AB1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[228*12+:12]), .o_data(A[228][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AB2_Mul0000000001(.i_data_1(c_plus_d[228][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[228][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AB3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[228*12+:12]), .o_data(C[228][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AB4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[484*12+:12]), .o_data(A[228][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AB5_Mul0000000001(.i_data_1(c_plus_d[228][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[228][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AB6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[484*12+:12]), .o_data(C[228][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AB7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[740*12+:12]), .o_data(A[228][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AB8_Mul0000000001(.i_data_1(c_plus_d[228][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[228][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AB9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[740*12+:12]), .o_data(C[228][2]), .i_clk(i_clk));
Mul0000000001  u_0000000ABA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[996*12+:12]), .o_data(A[228][3]), .i_clk(i_clk));
Mul0000000001  u_0000000ABB_Mul0000000001(.i_data_1(c_plus_d[228][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[228][3]), .i_clk(i_clk));
Mul0000000001  u_0000000ABC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[996*12+:12]), .o_data(C[228][3]), .i_clk(i_clk));
Mul0000000001  u_0000000ABD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[229*12+:12]), .o_data(A[229][0]), .i_clk(i_clk));
Mul0000000001  u_0000000ABE_Mul0000000001(.i_data_1(c_plus_d[229][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[229][0]), .i_clk(i_clk));
Mul0000000001  u_0000000ABF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[229*12+:12]), .o_data(C[229][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AC0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[485*12+:12]), .o_data(A[229][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AC1_Mul0000000001(.i_data_1(c_plus_d[229][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[229][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AC2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[485*12+:12]), .o_data(C[229][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AC3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[741*12+:12]), .o_data(A[229][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AC4_Mul0000000001(.i_data_1(c_plus_d[229][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[229][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AC5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[741*12+:12]), .o_data(C[229][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AC6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[997*12+:12]), .o_data(A[229][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AC7_Mul0000000001(.i_data_1(c_plus_d[229][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[229][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AC8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[997*12+:12]), .o_data(C[229][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AC9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[230*12+:12]), .o_data(A[230][0]), .i_clk(i_clk));
Mul0000000001  u_0000000ACA_Mul0000000001(.i_data_1(c_plus_d[230][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[230][0]), .i_clk(i_clk));
Mul0000000001  u_0000000ACB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[230*12+:12]), .o_data(C[230][0]), .i_clk(i_clk));
Mul0000000001  u_0000000ACC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[486*12+:12]), .o_data(A[230][1]), .i_clk(i_clk));
Mul0000000001  u_0000000ACD_Mul0000000001(.i_data_1(c_plus_d[230][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[230][1]), .i_clk(i_clk));
Mul0000000001  u_0000000ACE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[486*12+:12]), .o_data(C[230][1]), .i_clk(i_clk));
Mul0000000001  u_0000000ACF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[742*12+:12]), .o_data(A[230][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AD0_Mul0000000001(.i_data_1(c_plus_d[230][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[230][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AD1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[742*12+:12]), .o_data(C[230][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AD2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[998*12+:12]), .o_data(A[230][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AD3_Mul0000000001(.i_data_1(c_plus_d[230][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[230][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AD4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[998*12+:12]), .o_data(C[230][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AD5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[231*12+:12]), .o_data(A[231][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AD6_Mul0000000001(.i_data_1(c_plus_d[231][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[231][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AD7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[231*12+:12]), .o_data(C[231][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AD8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[487*12+:12]), .o_data(A[231][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AD9_Mul0000000001(.i_data_1(c_plus_d[231][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[231][1]), .i_clk(i_clk));
Mul0000000001  u_0000000ADA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[487*12+:12]), .o_data(C[231][1]), .i_clk(i_clk));
Mul0000000001  u_0000000ADB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[743*12+:12]), .o_data(A[231][2]), .i_clk(i_clk));
Mul0000000001  u_0000000ADC_Mul0000000001(.i_data_1(c_plus_d[231][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[231][2]), .i_clk(i_clk));
Mul0000000001  u_0000000ADD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[743*12+:12]), .o_data(C[231][2]), .i_clk(i_clk));
Mul0000000001  u_0000000ADE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[999*12+:12]), .o_data(A[231][3]), .i_clk(i_clk));
Mul0000000001  u_0000000ADF_Mul0000000001(.i_data_1(c_plus_d[231][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[231][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AE0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[999*12+:12]), .o_data(C[231][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AE1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[232*12+:12]), .o_data(A[232][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AE2_Mul0000000001(.i_data_1(c_plus_d[232][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[232][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AE3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[232*12+:12]), .o_data(C[232][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AE4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[488*12+:12]), .o_data(A[232][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AE5_Mul0000000001(.i_data_1(c_plus_d[232][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[232][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AE6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[488*12+:12]), .o_data(C[232][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AE7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[744*12+:12]), .o_data(A[232][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AE8_Mul0000000001(.i_data_1(c_plus_d[232][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[232][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AE9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[744*12+:12]), .o_data(C[232][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AEA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1000*12+:12]), .o_data(A[232][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AEB_Mul0000000001(.i_data_1(c_plus_d[232][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[232][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AEC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1000*12+:12]), .o_data(C[232][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AED_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[233*12+:12]), .o_data(A[233][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AEE_Mul0000000001(.i_data_1(c_plus_d[233][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[233][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AEF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[233*12+:12]), .o_data(C[233][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AF0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[489*12+:12]), .o_data(A[233][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AF1_Mul0000000001(.i_data_1(c_plus_d[233][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[233][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AF2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[489*12+:12]), .o_data(C[233][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AF3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[745*12+:12]), .o_data(A[233][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AF4_Mul0000000001(.i_data_1(c_plus_d[233][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[233][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AF5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[745*12+:12]), .o_data(C[233][2]), .i_clk(i_clk));
Mul0000000001  u_0000000AF6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1001*12+:12]), .o_data(A[233][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AF7_Mul0000000001(.i_data_1(c_plus_d[233][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[233][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AF8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1001*12+:12]), .o_data(C[233][3]), .i_clk(i_clk));
Mul0000000001  u_0000000AF9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[234*12+:12]), .o_data(A[234][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AFA_Mul0000000001(.i_data_1(c_plus_d[234][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[234][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AFB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[234*12+:12]), .o_data(C[234][0]), .i_clk(i_clk));
Mul0000000001  u_0000000AFC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[490*12+:12]), .o_data(A[234][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AFD_Mul0000000001(.i_data_1(c_plus_d[234][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[234][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AFE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[490*12+:12]), .o_data(C[234][1]), .i_clk(i_clk));
Mul0000000001  u_0000000AFF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[746*12+:12]), .o_data(A[234][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B00_Mul0000000001(.i_data_1(c_plus_d[234][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[234][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B01_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[746*12+:12]), .o_data(C[234][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B02_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1002*12+:12]), .o_data(A[234][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B03_Mul0000000001(.i_data_1(c_plus_d[234][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[234][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B04_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1002*12+:12]), .o_data(C[234][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B05_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[235*12+:12]), .o_data(A[235][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B06_Mul0000000001(.i_data_1(c_plus_d[235][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[235][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B07_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[235*12+:12]), .o_data(C[235][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B08_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[491*12+:12]), .o_data(A[235][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B09_Mul0000000001(.i_data_1(c_plus_d[235][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[235][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B0A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[491*12+:12]), .o_data(C[235][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B0B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[747*12+:12]), .o_data(A[235][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B0C_Mul0000000001(.i_data_1(c_plus_d[235][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[235][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B0D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[747*12+:12]), .o_data(C[235][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B0E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1003*12+:12]), .o_data(A[235][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B0F_Mul0000000001(.i_data_1(c_plus_d[235][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[235][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B10_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1003*12+:12]), .o_data(C[235][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B11_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[236*12+:12]), .o_data(A[236][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B12_Mul0000000001(.i_data_1(c_plus_d[236][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[236][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B13_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[236*12+:12]), .o_data(C[236][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B14_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[492*12+:12]), .o_data(A[236][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B15_Mul0000000001(.i_data_1(c_plus_d[236][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[236][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B16_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[492*12+:12]), .o_data(C[236][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B17_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[748*12+:12]), .o_data(A[236][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B18_Mul0000000001(.i_data_1(c_plus_d[236][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[236][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B19_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[748*12+:12]), .o_data(C[236][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B1A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1004*12+:12]), .o_data(A[236][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B1B_Mul0000000001(.i_data_1(c_plus_d[236][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[236][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B1C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1004*12+:12]), .o_data(C[236][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B1D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[237*12+:12]), .o_data(A[237][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B1E_Mul0000000001(.i_data_1(c_plus_d[237][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[237][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B1F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[237*12+:12]), .o_data(C[237][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B20_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[493*12+:12]), .o_data(A[237][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B21_Mul0000000001(.i_data_1(c_plus_d[237][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[237][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B22_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[493*12+:12]), .o_data(C[237][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B23_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[749*12+:12]), .o_data(A[237][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B24_Mul0000000001(.i_data_1(c_plus_d[237][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[237][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B25_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[749*12+:12]), .o_data(C[237][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B26_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1005*12+:12]), .o_data(A[237][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B27_Mul0000000001(.i_data_1(c_plus_d[237][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[237][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B28_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1005*12+:12]), .o_data(C[237][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B29_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[238*12+:12]), .o_data(A[238][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B2A_Mul0000000001(.i_data_1(c_plus_d[238][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[238][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B2B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[238*12+:12]), .o_data(C[238][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B2C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[494*12+:12]), .o_data(A[238][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B2D_Mul0000000001(.i_data_1(c_plus_d[238][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[238][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B2E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[494*12+:12]), .o_data(C[238][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B2F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[750*12+:12]), .o_data(A[238][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B30_Mul0000000001(.i_data_1(c_plus_d[238][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[238][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B31_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[750*12+:12]), .o_data(C[238][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B32_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1006*12+:12]), .o_data(A[238][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B33_Mul0000000001(.i_data_1(c_plus_d[238][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[238][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B34_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1006*12+:12]), .o_data(C[238][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B35_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[239*12+:12]), .o_data(A[239][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B36_Mul0000000001(.i_data_1(c_plus_d[239][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[239][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B37_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[239*12+:12]), .o_data(C[239][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B38_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[495*12+:12]), .o_data(A[239][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B39_Mul0000000001(.i_data_1(c_plus_d[239][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[239][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B3A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[495*12+:12]), .o_data(C[239][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B3B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[751*12+:12]), .o_data(A[239][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B3C_Mul0000000001(.i_data_1(c_plus_d[239][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[239][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B3D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[751*12+:12]), .o_data(C[239][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B3E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1007*12+:12]), .o_data(A[239][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B3F_Mul0000000001(.i_data_1(c_plus_d[239][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[239][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B40_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1007*12+:12]), .o_data(C[239][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B41_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[240*12+:12]), .o_data(A[240][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B42_Mul0000000001(.i_data_1(c_plus_d[240][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[240][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B43_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[240*12+:12]), .o_data(C[240][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B44_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[496*12+:12]), .o_data(A[240][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B45_Mul0000000001(.i_data_1(c_plus_d[240][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[240][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B46_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[496*12+:12]), .o_data(C[240][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B47_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[752*12+:12]), .o_data(A[240][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B48_Mul0000000001(.i_data_1(c_plus_d[240][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[240][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B49_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[752*12+:12]), .o_data(C[240][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B4A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1008*12+:12]), .o_data(A[240][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B4B_Mul0000000001(.i_data_1(c_plus_d[240][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[240][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B4C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1008*12+:12]), .o_data(C[240][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B4D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[241*12+:12]), .o_data(A[241][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B4E_Mul0000000001(.i_data_1(c_plus_d[241][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[241][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B4F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[241*12+:12]), .o_data(C[241][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B50_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[497*12+:12]), .o_data(A[241][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B51_Mul0000000001(.i_data_1(c_plus_d[241][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[241][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B52_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[497*12+:12]), .o_data(C[241][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B53_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[753*12+:12]), .o_data(A[241][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B54_Mul0000000001(.i_data_1(c_plus_d[241][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[241][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B55_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[753*12+:12]), .o_data(C[241][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B56_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1009*12+:12]), .o_data(A[241][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B57_Mul0000000001(.i_data_1(c_plus_d[241][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[241][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B58_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1009*12+:12]), .o_data(C[241][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B59_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[242*12+:12]), .o_data(A[242][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B5A_Mul0000000001(.i_data_1(c_plus_d[242][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[242][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B5B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[242*12+:12]), .o_data(C[242][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B5C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[498*12+:12]), .o_data(A[242][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B5D_Mul0000000001(.i_data_1(c_plus_d[242][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[242][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B5E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[498*12+:12]), .o_data(C[242][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B5F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[754*12+:12]), .o_data(A[242][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B60_Mul0000000001(.i_data_1(c_plus_d[242][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[242][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B61_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[754*12+:12]), .o_data(C[242][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B62_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1010*12+:12]), .o_data(A[242][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B63_Mul0000000001(.i_data_1(c_plus_d[242][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[242][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B64_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1010*12+:12]), .o_data(C[242][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B65_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[243*12+:12]), .o_data(A[243][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B66_Mul0000000001(.i_data_1(c_plus_d[243][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[243][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B67_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[243*12+:12]), .o_data(C[243][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B68_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[499*12+:12]), .o_data(A[243][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B69_Mul0000000001(.i_data_1(c_plus_d[243][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[243][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B6A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[499*12+:12]), .o_data(C[243][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B6B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[755*12+:12]), .o_data(A[243][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B6C_Mul0000000001(.i_data_1(c_plus_d[243][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[243][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B6D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[755*12+:12]), .o_data(C[243][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B6E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1011*12+:12]), .o_data(A[243][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B6F_Mul0000000001(.i_data_1(c_plus_d[243][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[243][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B70_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1011*12+:12]), .o_data(C[243][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B71_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[244*12+:12]), .o_data(A[244][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B72_Mul0000000001(.i_data_1(c_plus_d[244][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[244][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B73_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[244*12+:12]), .o_data(C[244][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B74_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[500*12+:12]), .o_data(A[244][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B75_Mul0000000001(.i_data_1(c_plus_d[244][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[244][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B76_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[500*12+:12]), .o_data(C[244][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B77_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[756*12+:12]), .o_data(A[244][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B78_Mul0000000001(.i_data_1(c_plus_d[244][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[244][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B79_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[756*12+:12]), .o_data(C[244][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B7A_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1012*12+:12]), .o_data(A[244][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B7B_Mul0000000001(.i_data_1(c_plus_d[244][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[244][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B7C_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1012*12+:12]), .o_data(C[244][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B7D_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[245*12+:12]), .o_data(A[245][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B7E_Mul0000000001(.i_data_1(c_plus_d[245][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[245][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B7F_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[245*12+:12]), .o_data(C[245][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B80_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[501*12+:12]), .o_data(A[245][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B81_Mul0000000001(.i_data_1(c_plus_d[245][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[245][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B82_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[501*12+:12]), .o_data(C[245][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B83_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[757*12+:12]), .o_data(A[245][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B84_Mul0000000001(.i_data_1(c_plus_d[245][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[245][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B85_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[757*12+:12]), .o_data(C[245][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B86_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1013*12+:12]), .o_data(A[245][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B87_Mul0000000001(.i_data_1(c_plus_d[245][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[245][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B88_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1013*12+:12]), .o_data(C[245][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B89_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[246*12+:12]), .o_data(A[246][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B8A_Mul0000000001(.i_data_1(c_plus_d[246][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[246][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B8B_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[246*12+:12]), .o_data(C[246][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B8C_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[502*12+:12]), .o_data(A[246][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B8D_Mul0000000001(.i_data_1(c_plus_d[246][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[246][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B8E_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[502*12+:12]), .o_data(C[246][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B8F_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[758*12+:12]), .o_data(A[246][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B90_Mul0000000001(.i_data_1(c_plus_d[246][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[246][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B91_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[758*12+:12]), .o_data(C[246][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B92_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1014*12+:12]), .o_data(A[246][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B93_Mul0000000001(.i_data_1(c_plus_d[246][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[246][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B94_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1014*12+:12]), .o_data(C[246][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B95_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[247*12+:12]), .o_data(A[247][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B96_Mul0000000001(.i_data_1(c_plus_d[247][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[247][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B97_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[247*12+:12]), .o_data(C[247][0]), .i_clk(i_clk));
Mul0000000001  u_0000000B98_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[503*12+:12]), .o_data(A[247][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B99_Mul0000000001(.i_data_1(c_plus_d[247][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[247][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B9A_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[503*12+:12]), .o_data(C[247][1]), .i_clk(i_clk));
Mul0000000001  u_0000000B9B_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[759*12+:12]), .o_data(A[247][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B9C_Mul0000000001(.i_data_1(c_plus_d[247][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[247][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B9D_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[759*12+:12]), .o_data(C[247][2]), .i_clk(i_clk));
Mul0000000001  u_0000000B9E_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1015*12+:12]), .o_data(A[247][3]), .i_clk(i_clk));
Mul0000000001  u_0000000B9F_Mul0000000001(.i_data_1(c_plus_d[247][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[247][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BA0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1015*12+:12]), .o_data(C[247][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BA1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[248*12+:12]), .o_data(A[248][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BA2_Mul0000000001(.i_data_1(c_plus_d[248][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[248][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BA3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[248*12+:12]), .o_data(C[248][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BA4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[504*12+:12]), .o_data(A[248][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BA5_Mul0000000001(.i_data_1(c_plus_d[248][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[248][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BA6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[504*12+:12]), .o_data(C[248][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BA7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[760*12+:12]), .o_data(A[248][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BA8_Mul0000000001(.i_data_1(c_plus_d[248][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[248][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BA9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[760*12+:12]), .o_data(C[248][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BAA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1016*12+:12]), .o_data(A[248][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BAB_Mul0000000001(.i_data_1(c_plus_d[248][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[248][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BAC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1016*12+:12]), .o_data(C[248][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BAD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[249*12+:12]), .o_data(A[249][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BAE_Mul0000000001(.i_data_1(c_plus_d[249][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[249][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BAF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[249*12+:12]), .o_data(C[249][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BB0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[505*12+:12]), .o_data(A[249][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BB1_Mul0000000001(.i_data_1(c_plus_d[249][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[249][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BB2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[505*12+:12]), .o_data(C[249][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BB3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[761*12+:12]), .o_data(A[249][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BB4_Mul0000000001(.i_data_1(c_plus_d[249][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[249][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BB5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[761*12+:12]), .o_data(C[249][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BB6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1017*12+:12]), .o_data(A[249][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BB7_Mul0000000001(.i_data_1(c_plus_d[249][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[249][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BB8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1017*12+:12]), .o_data(C[249][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BB9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[250*12+:12]), .o_data(A[250][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BBA_Mul0000000001(.i_data_1(c_plus_d[250][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[250][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BBB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[250*12+:12]), .o_data(C[250][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BBC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[506*12+:12]), .o_data(A[250][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BBD_Mul0000000001(.i_data_1(c_plus_d[250][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[250][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BBE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[506*12+:12]), .o_data(C[250][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BBF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[762*12+:12]), .o_data(A[250][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BC0_Mul0000000001(.i_data_1(c_plus_d[250][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[250][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BC1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[762*12+:12]), .o_data(C[250][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BC2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1018*12+:12]), .o_data(A[250][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BC3_Mul0000000001(.i_data_1(c_plus_d[250][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[250][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BC4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1018*12+:12]), .o_data(C[250][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BC5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[251*12+:12]), .o_data(A[251][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BC6_Mul0000000001(.i_data_1(c_plus_d[251][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[251][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BC7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[251*12+:12]), .o_data(C[251][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BC8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[507*12+:12]), .o_data(A[251][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BC9_Mul0000000001(.i_data_1(c_plus_d[251][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[251][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BCA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[507*12+:12]), .o_data(C[251][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BCB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[763*12+:12]), .o_data(A[251][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BCC_Mul0000000001(.i_data_1(c_plus_d[251][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[251][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BCD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[763*12+:12]), .o_data(C[251][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BCE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1019*12+:12]), .o_data(A[251][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BCF_Mul0000000001(.i_data_1(c_plus_d[251][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[251][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BD0_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1019*12+:12]), .o_data(C[251][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BD1_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[252*12+:12]), .o_data(A[252][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BD2_Mul0000000001(.i_data_1(c_plus_d[252][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[252][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BD3_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[252*12+:12]), .o_data(C[252][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BD4_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[508*12+:12]), .o_data(A[252][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BD5_Mul0000000001(.i_data_1(c_plus_d[252][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[252][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BD6_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[508*12+:12]), .o_data(C[252][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BD7_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[764*12+:12]), .o_data(A[252][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BD8_Mul0000000001(.i_data_1(c_plus_d[252][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[252][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BD9_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[764*12+:12]), .o_data(C[252][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BDA_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1020*12+:12]), .o_data(A[252][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BDB_Mul0000000001(.i_data_1(c_plus_d[252][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[252][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BDC_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1020*12+:12]), .o_data(C[252][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BDD_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[253*12+:12]), .o_data(A[253][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BDE_Mul0000000001(.i_data_1(c_plus_d[253][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[253][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BDF_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[253*12+:12]), .o_data(C[253][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BE0_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[509*12+:12]), .o_data(A[253][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BE1_Mul0000000001(.i_data_1(c_plus_d[253][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[253][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BE2_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[509*12+:12]), .o_data(C[253][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BE3_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[765*12+:12]), .o_data(A[253][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BE4_Mul0000000001(.i_data_1(c_plus_d[253][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[253][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BE5_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[765*12+:12]), .o_data(C[253][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BE6_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1021*12+:12]), .o_data(A[253][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BE7_Mul0000000001(.i_data_1(c_plus_d[253][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[253][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BE8_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1021*12+:12]), .o_data(C[253][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BE9_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[254*12+:12]), .o_data(A[254][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BEA_Mul0000000001(.i_data_1(c_plus_d[254][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[254][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BEB_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[254*12+:12]), .o_data(C[254][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BEC_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[510*12+:12]), .o_data(A[254][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BED_Mul0000000001(.i_data_1(c_plus_d[254][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[254][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BEE_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[510*12+:12]), .o_data(C[254][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BEF_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[766*12+:12]), .o_data(A[254][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BF0_Mul0000000001(.i_data_1(c_plus_d[254][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[254][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BF1_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[766*12+:12]), .o_data(C[254][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BF2_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1022*12+:12]), .o_data(A[254][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BF3_Mul0000000001(.i_data_1(c_plus_d[254][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[254][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BF4_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1022*12+:12]), .o_data(C[254][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BF5_Mul0000000001(.i_data_1(a_plus_b[0]), .i_data_2(matrix_r_d[255*12+:12]), .o_data(A[255][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BF6_Mul0000000001(.i_data_1(c_plus_d[255][0]), .i_data_2(vector_i_d[0*12+:12]), .o_data(B[255][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BF7_Mul0000000001(.i_data_1(b_minus_a[0]), .i_data_2(matrix_i_d[255*12+:12]), .o_data(C[255][0]), .i_clk(i_clk));
Mul0000000001  u_0000000BF8_Mul0000000001(.i_data_1(a_plus_b[1]), .i_data_2(matrix_r_d[511*12+:12]), .o_data(A[255][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BF9_Mul0000000001(.i_data_1(c_plus_d[255][1]), .i_data_2(vector_i_d[1*12+:12]), .o_data(B[255][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BFA_Mul0000000001(.i_data_1(b_minus_a[1]), .i_data_2(matrix_i_d[511*12+:12]), .o_data(C[255][1]), .i_clk(i_clk));
Mul0000000001  u_0000000BFB_Mul0000000001(.i_data_1(a_plus_b[2]), .i_data_2(matrix_r_d[767*12+:12]), .o_data(A[255][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BFC_Mul0000000001(.i_data_1(c_plus_d[255][2]), .i_data_2(vector_i_d[2*12+:12]), .o_data(B[255][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BFD_Mul0000000001(.i_data_1(b_minus_a[2]), .i_data_2(matrix_i_d[767*12+:12]), .o_data(C[255][2]), .i_clk(i_clk));
Mul0000000001  u_0000000BFE_Mul0000000001(.i_data_1(a_plus_b[3]), .i_data_2(matrix_r_d[1023*12+:12]), .o_data(A[255][3]), .i_clk(i_clk));
Mul0000000001  u_0000000BFF_Mul0000000001(.i_data_1(c_plus_d[255][3]), .i_data_2(vector_i_d[3*12+:12]), .o_data(B[255][3]), .i_clk(i_clk));
Mul0000000001  u_0000000C00_Mul0000000001(.i_data_1(b_minus_a[3]), .i_data_2(matrix_i_d[1023*12+:12]), .o_data(C[255][3]), .i_clk(i_clk));
 // Layer 3: Subtraction
 wire [12-1:0] mult_result_r [0:256-1][0:4-1];
 wire [12-1:0] mult_result_i [0:256-1][0:4-1];
Sub0000000002  u_0000000001_Sub0000000002(.i_data_1(A[0][0]), .i_data_2(B[0][0]), .o_data(mult_result_r[0][0]), .i_clk(i_clk));
Sub0000000002  u_0000000002_Sub0000000002(.i_data_1(B[0][0]), .i_data_2(C[0][0]), .o_data(mult_result_i[0][0]), .i_clk(i_clk));
Sub0000000002  u_0000000003_Sub0000000002(.i_data_1(A[0][1]), .i_data_2(B[0][1]), .o_data(mult_result_r[0][1]), .i_clk(i_clk));
Sub0000000002  u_0000000004_Sub0000000002(.i_data_1(B[0][1]), .i_data_2(C[0][1]), .o_data(mult_result_i[0][1]), .i_clk(i_clk));
Sub0000000002  u_0000000005_Sub0000000002(.i_data_1(A[0][2]), .i_data_2(B[0][2]), .o_data(mult_result_r[0][2]), .i_clk(i_clk));
Sub0000000002  u_0000000006_Sub0000000002(.i_data_1(B[0][2]), .i_data_2(C[0][2]), .o_data(mult_result_i[0][2]), .i_clk(i_clk));
Sub0000000002  u_0000000007_Sub0000000002(.i_data_1(A[0][3]), .i_data_2(B[0][3]), .o_data(mult_result_r[0][3]), .i_clk(i_clk));
Sub0000000002  u_0000000008_Sub0000000002(.i_data_1(B[0][3]), .i_data_2(C[0][3]), .o_data(mult_result_i[0][3]), .i_clk(i_clk));
Sub0000000002  u_0000000009_Sub0000000002(.i_data_1(A[1][0]), .i_data_2(B[1][0]), .o_data(mult_result_r[1][0]), .i_clk(i_clk));
Sub0000000002  u_000000000A_Sub0000000002(.i_data_1(B[1][0]), .i_data_2(C[1][0]), .o_data(mult_result_i[1][0]), .i_clk(i_clk));
Sub0000000002  u_000000000B_Sub0000000002(.i_data_1(A[1][1]), .i_data_2(B[1][1]), .o_data(mult_result_r[1][1]), .i_clk(i_clk));
Sub0000000002  u_000000000C_Sub0000000002(.i_data_1(B[1][1]), .i_data_2(C[1][1]), .o_data(mult_result_i[1][1]), .i_clk(i_clk));
Sub0000000002  u_000000000D_Sub0000000002(.i_data_1(A[1][2]), .i_data_2(B[1][2]), .o_data(mult_result_r[1][2]), .i_clk(i_clk));
Sub0000000002  u_000000000E_Sub0000000002(.i_data_1(B[1][2]), .i_data_2(C[1][2]), .o_data(mult_result_i[1][2]), .i_clk(i_clk));
Sub0000000002  u_000000000F_Sub0000000002(.i_data_1(A[1][3]), .i_data_2(B[1][3]), .o_data(mult_result_r[1][3]), .i_clk(i_clk));
Sub0000000002  u_0000000010_Sub0000000002(.i_data_1(B[1][3]), .i_data_2(C[1][3]), .o_data(mult_result_i[1][3]), .i_clk(i_clk));
Sub0000000002  u_0000000011_Sub0000000002(.i_data_1(A[2][0]), .i_data_2(B[2][0]), .o_data(mult_result_r[2][0]), .i_clk(i_clk));
Sub0000000002  u_0000000012_Sub0000000002(.i_data_1(B[2][0]), .i_data_2(C[2][0]), .o_data(mult_result_i[2][0]), .i_clk(i_clk));
Sub0000000002  u_0000000013_Sub0000000002(.i_data_1(A[2][1]), .i_data_2(B[2][1]), .o_data(mult_result_r[2][1]), .i_clk(i_clk));
Sub0000000002  u_0000000014_Sub0000000002(.i_data_1(B[2][1]), .i_data_2(C[2][1]), .o_data(mult_result_i[2][1]), .i_clk(i_clk));
Sub0000000002  u_0000000015_Sub0000000002(.i_data_1(A[2][2]), .i_data_2(B[2][2]), .o_data(mult_result_r[2][2]), .i_clk(i_clk));
Sub0000000002  u_0000000016_Sub0000000002(.i_data_1(B[2][2]), .i_data_2(C[2][2]), .o_data(mult_result_i[2][2]), .i_clk(i_clk));
Sub0000000002  u_0000000017_Sub0000000002(.i_data_1(A[2][3]), .i_data_2(B[2][3]), .o_data(mult_result_r[2][3]), .i_clk(i_clk));
Sub0000000002  u_0000000018_Sub0000000002(.i_data_1(B[2][3]), .i_data_2(C[2][3]), .o_data(mult_result_i[2][3]), .i_clk(i_clk));
Sub0000000002  u_0000000019_Sub0000000002(.i_data_1(A[3][0]), .i_data_2(B[3][0]), .o_data(mult_result_r[3][0]), .i_clk(i_clk));
Sub0000000002  u_000000001A_Sub0000000002(.i_data_1(B[3][0]), .i_data_2(C[3][0]), .o_data(mult_result_i[3][0]), .i_clk(i_clk));
Sub0000000002  u_000000001B_Sub0000000002(.i_data_1(A[3][1]), .i_data_2(B[3][1]), .o_data(mult_result_r[3][1]), .i_clk(i_clk));
Sub0000000002  u_000000001C_Sub0000000002(.i_data_1(B[3][1]), .i_data_2(C[3][1]), .o_data(mult_result_i[3][1]), .i_clk(i_clk));
Sub0000000002  u_000000001D_Sub0000000002(.i_data_1(A[3][2]), .i_data_2(B[3][2]), .o_data(mult_result_r[3][2]), .i_clk(i_clk));
Sub0000000002  u_000000001E_Sub0000000002(.i_data_1(B[3][2]), .i_data_2(C[3][2]), .o_data(mult_result_i[3][2]), .i_clk(i_clk));
Sub0000000002  u_000000001F_Sub0000000002(.i_data_1(A[3][3]), .i_data_2(B[3][3]), .o_data(mult_result_r[3][3]), .i_clk(i_clk));
Sub0000000002  u_0000000020_Sub0000000002(.i_data_1(B[3][3]), .i_data_2(C[3][3]), .o_data(mult_result_i[3][3]), .i_clk(i_clk));
Sub0000000002  u_0000000021_Sub0000000002(.i_data_1(A[4][0]), .i_data_2(B[4][0]), .o_data(mult_result_r[4][0]), .i_clk(i_clk));
Sub0000000002  u_0000000022_Sub0000000002(.i_data_1(B[4][0]), .i_data_2(C[4][0]), .o_data(mult_result_i[4][0]), .i_clk(i_clk));
Sub0000000002  u_0000000023_Sub0000000002(.i_data_1(A[4][1]), .i_data_2(B[4][1]), .o_data(mult_result_r[4][1]), .i_clk(i_clk));
Sub0000000002  u_0000000024_Sub0000000002(.i_data_1(B[4][1]), .i_data_2(C[4][1]), .o_data(mult_result_i[4][1]), .i_clk(i_clk));
Sub0000000002  u_0000000025_Sub0000000002(.i_data_1(A[4][2]), .i_data_2(B[4][2]), .o_data(mult_result_r[4][2]), .i_clk(i_clk));
Sub0000000002  u_0000000026_Sub0000000002(.i_data_1(B[4][2]), .i_data_2(C[4][2]), .o_data(mult_result_i[4][2]), .i_clk(i_clk));
Sub0000000002  u_0000000027_Sub0000000002(.i_data_1(A[4][3]), .i_data_2(B[4][3]), .o_data(mult_result_r[4][3]), .i_clk(i_clk));
Sub0000000002  u_0000000028_Sub0000000002(.i_data_1(B[4][3]), .i_data_2(C[4][3]), .o_data(mult_result_i[4][3]), .i_clk(i_clk));
Sub0000000002  u_0000000029_Sub0000000002(.i_data_1(A[5][0]), .i_data_2(B[5][0]), .o_data(mult_result_r[5][0]), .i_clk(i_clk));
Sub0000000002  u_000000002A_Sub0000000002(.i_data_1(B[5][0]), .i_data_2(C[5][0]), .o_data(mult_result_i[5][0]), .i_clk(i_clk));
Sub0000000002  u_000000002B_Sub0000000002(.i_data_1(A[5][1]), .i_data_2(B[5][1]), .o_data(mult_result_r[5][1]), .i_clk(i_clk));
Sub0000000002  u_000000002C_Sub0000000002(.i_data_1(B[5][1]), .i_data_2(C[5][1]), .o_data(mult_result_i[5][1]), .i_clk(i_clk));
Sub0000000002  u_000000002D_Sub0000000002(.i_data_1(A[5][2]), .i_data_2(B[5][2]), .o_data(mult_result_r[5][2]), .i_clk(i_clk));
Sub0000000002  u_000000002E_Sub0000000002(.i_data_1(B[5][2]), .i_data_2(C[5][2]), .o_data(mult_result_i[5][2]), .i_clk(i_clk));
Sub0000000002  u_000000002F_Sub0000000002(.i_data_1(A[5][3]), .i_data_2(B[5][3]), .o_data(mult_result_r[5][3]), .i_clk(i_clk));
Sub0000000002  u_0000000030_Sub0000000002(.i_data_1(B[5][3]), .i_data_2(C[5][3]), .o_data(mult_result_i[5][3]), .i_clk(i_clk));
Sub0000000002  u_0000000031_Sub0000000002(.i_data_1(A[6][0]), .i_data_2(B[6][0]), .o_data(mult_result_r[6][0]), .i_clk(i_clk));
Sub0000000002  u_0000000032_Sub0000000002(.i_data_1(B[6][0]), .i_data_2(C[6][0]), .o_data(mult_result_i[6][0]), .i_clk(i_clk));
Sub0000000002  u_0000000033_Sub0000000002(.i_data_1(A[6][1]), .i_data_2(B[6][1]), .o_data(mult_result_r[6][1]), .i_clk(i_clk));
Sub0000000002  u_0000000034_Sub0000000002(.i_data_1(B[6][1]), .i_data_2(C[6][1]), .o_data(mult_result_i[6][1]), .i_clk(i_clk));
Sub0000000002  u_0000000035_Sub0000000002(.i_data_1(A[6][2]), .i_data_2(B[6][2]), .o_data(mult_result_r[6][2]), .i_clk(i_clk));
Sub0000000002  u_0000000036_Sub0000000002(.i_data_1(B[6][2]), .i_data_2(C[6][2]), .o_data(mult_result_i[6][2]), .i_clk(i_clk));
Sub0000000002  u_0000000037_Sub0000000002(.i_data_1(A[6][3]), .i_data_2(B[6][3]), .o_data(mult_result_r[6][3]), .i_clk(i_clk));
Sub0000000002  u_0000000038_Sub0000000002(.i_data_1(B[6][3]), .i_data_2(C[6][3]), .o_data(mult_result_i[6][3]), .i_clk(i_clk));
Sub0000000002  u_0000000039_Sub0000000002(.i_data_1(A[7][0]), .i_data_2(B[7][0]), .o_data(mult_result_r[7][0]), .i_clk(i_clk));
Sub0000000002  u_000000003A_Sub0000000002(.i_data_1(B[7][0]), .i_data_2(C[7][0]), .o_data(mult_result_i[7][0]), .i_clk(i_clk));
Sub0000000002  u_000000003B_Sub0000000002(.i_data_1(A[7][1]), .i_data_2(B[7][1]), .o_data(mult_result_r[7][1]), .i_clk(i_clk));
Sub0000000002  u_000000003C_Sub0000000002(.i_data_1(B[7][1]), .i_data_2(C[7][1]), .o_data(mult_result_i[7][1]), .i_clk(i_clk));
Sub0000000002  u_000000003D_Sub0000000002(.i_data_1(A[7][2]), .i_data_2(B[7][2]), .o_data(mult_result_r[7][2]), .i_clk(i_clk));
Sub0000000002  u_000000003E_Sub0000000002(.i_data_1(B[7][2]), .i_data_2(C[7][2]), .o_data(mult_result_i[7][2]), .i_clk(i_clk));
Sub0000000002  u_000000003F_Sub0000000002(.i_data_1(A[7][3]), .i_data_2(B[7][3]), .o_data(mult_result_r[7][3]), .i_clk(i_clk));
Sub0000000002  u_0000000040_Sub0000000002(.i_data_1(B[7][3]), .i_data_2(C[7][3]), .o_data(mult_result_i[7][3]), .i_clk(i_clk));
Sub0000000002  u_0000000041_Sub0000000002(.i_data_1(A[8][0]), .i_data_2(B[8][0]), .o_data(mult_result_r[8][0]), .i_clk(i_clk));
Sub0000000002  u_0000000042_Sub0000000002(.i_data_1(B[8][0]), .i_data_2(C[8][0]), .o_data(mult_result_i[8][0]), .i_clk(i_clk));
Sub0000000002  u_0000000043_Sub0000000002(.i_data_1(A[8][1]), .i_data_2(B[8][1]), .o_data(mult_result_r[8][1]), .i_clk(i_clk));
Sub0000000002  u_0000000044_Sub0000000002(.i_data_1(B[8][1]), .i_data_2(C[8][1]), .o_data(mult_result_i[8][1]), .i_clk(i_clk));
Sub0000000002  u_0000000045_Sub0000000002(.i_data_1(A[8][2]), .i_data_2(B[8][2]), .o_data(mult_result_r[8][2]), .i_clk(i_clk));
Sub0000000002  u_0000000046_Sub0000000002(.i_data_1(B[8][2]), .i_data_2(C[8][2]), .o_data(mult_result_i[8][2]), .i_clk(i_clk));
Sub0000000002  u_0000000047_Sub0000000002(.i_data_1(A[8][3]), .i_data_2(B[8][3]), .o_data(mult_result_r[8][3]), .i_clk(i_clk));
Sub0000000002  u_0000000048_Sub0000000002(.i_data_1(B[8][3]), .i_data_2(C[8][3]), .o_data(mult_result_i[8][3]), .i_clk(i_clk));
Sub0000000002  u_0000000049_Sub0000000002(.i_data_1(A[9][0]), .i_data_2(B[9][0]), .o_data(mult_result_r[9][0]), .i_clk(i_clk));
Sub0000000002  u_000000004A_Sub0000000002(.i_data_1(B[9][0]), .i_data_2(C[9][0]), .o_data(mult_result_i[9][0]), .i_clk(i_clk));
Sub0000000002  u_000000004B_Sub0000000002(.i_data_1(A[9][1]), .i_data_2(B[9][1]), .o_data(mult_result_r[9][1]), .i_clk(i_clk));
Sub0000000002  u_000000004C_Sub0000000002(.i_data_1(B[9][1]), .i_data_2(C[9][1]), .o_data(mult_result_i[9][1]), .i_clk(i_clk));
Sub0000000002  u_000000004D_Sub0000000002(.i_data_1(A[9][2]), .i_data_2(B[9][2]), .o_data(mult_result_r[9][2]), .i_clk(i_clk));
Sub0000000002  u_000000004E_Sub0000000002(.i_data_1(B[9][2]), .i_data_2(C[9][2]), .o_data(mult_result_i[9][2]), .i_clk(i_clk));
Sub0000000002  u_000000004F_Sub0000000002(.i_data_1(A[9][3]), .i_data_2(B[9][3]), .o_data(mult_result_r[9][3]), .i_clk(i_clk));
Sub0000000002  u_0000000050_Sub0000000002(.i_data_1(B[9][3]), .i_data_2(C[9][3]), .o_data(mult_result_i[9][3]), .i_clk(i_clk));
Sub0000000002  u_0000000051_Sub0000000002(.i_data_1(A[10][0]), .i_data_2(B[10][0]), .o_data(mult_result_r[10][0]), .i_clk(i_clk));
Sub0000000002  u_0000000052_Sub0000000002(.i_data_1(B[10][0]), .i_data_2(C[10][0]), .o_data(mult_result_i[10][0]), .i_clk(i_clk));
Sub0000000002  u_0000000053_Sub0000000002(.i_data_1(A[10][1]), .i_data_2(B[10][1]), .o_data(mult_result_r[10][1]), .i_clk(i_clk));
Sub0000000002  u_0000000054_Sub0000000002(.i_data_1(B[10][1]), .i_data_2(C[10][1]), .o_data(mult_result_i[10][1]), .i_clk(i_clk));
Sub0000000002  u_0000000055_Sub0000000002(.i_data_1(A[10][2]), .i_data_2(B[10][2]), .o_data(mult_result_r[10][2]), .i_clk(i_clk));
Sub0000000002  u_0000000056_Sub0000000002(.i_data_1(B[10][2]), .i_data_2(C[10][2]), .o_data(mult_result_i[10][2]), .i_clk(i_clk));
Sub0000000002  u_0000000057_Sub0000000002(.i_data_1(A[10][3]), .i_data_2(B[10][3]), .o_data(mult_result_r[10][3]), .i_clk(i_clk));
Sub0000000002  u_0000000058_Sub0000000002(.i_data_1(B[10][3]), .i_data_2(C[10][3]), .o_data(mult_result_i[10][3]), .i_clk(i_clk));
Sub0000000002  u_0000000059_Sub0000000002(.i_data_1(A[11][0]), .i_data_2(B[11][0]), .o_data(mult_result_r[11][0]), .i_clk(i_clk));
Sub0000000002  u_000000005A_Sub0000000002(.i_data_1(B[11][0]), .i_data_2(C[11][0]), .o_data(mult_result_i[11][0]), .i_clk(i_clk));
Sub0000000002  u_000000005B_Sub0000000002(.i_data_1(A[11][1]), .i_data_2(B[11][1]), .o_data(mult_result_r[11][1]), .i_clk(i_clk));
Sub0000000002  u_000000005C_Sub0000000002(.i_data_1(B[11][1]), .i_data_2(C[11][1]), .o_data(mult_result_i[11][1]), .i_clk(i_clk));
Sub0000000002  u_000000005D_Sub0000000002(.i_data_1(A[11][2]), .i_data_2(B[11][2]), .o_data(mult_result_r[11][2]), .i_clk(i_clk));
Sub0000000002  u_000000005E_Sub0000000002(.i_data_1(B[11][2]), .i_data_2(C[11][2]), .o_data(mult_result_i[11][2]), .i_clk(i_clk));
Sub0000000002  u_000000005F_Sub0000000002(.i_data_1(A[11][3]), .i_data_2(B[11][3]), .o_data(mult_result_r[11][3]), .i_clk(i_clk));
Sub0000000002  u_0000000060_Sub0000000002(.i_data_1(B[11][3]), .i_data_2(C[11][3]), .o_data(mult_result_i[11][3]), .i_clk(i_clk));
Sub0000000002  u_0000000061_Sub0000000002(.i_data_1(A[12][0]), .i_data_2(B[12][0]), .o_data(mult_result_r[12][0]), .i_clk(i_clk));
Sub0000000002  u_0000000062_Sub0000000002(.i_data_1(B[12][0]), .i_data_2(C[12][0]), .o_data(mult_result_i[12][0]), .i_clk(i_clk));
Sub0000000002  u_0000000063_Sub0000000002(.i_data_1(A[12][1]), .i_data_2(B[12][1]), .o_data(mult_result_r[12][1]), .i_clk(i_clk));
Sub0000000002  u_0000000064_Sub0000000002(.i_data_1(B[12][1]), .i_data_2(C[12][1]), .o_data(mult_result_i[12][1]), .i_clk(i_clk));
Sub0000000002  u_0000000065_Sub0000000002(.i_data_1(A[12][2]), .i_data_2(B[12][2]), .o_data(mult_result_r[12][2]), .i_clk(i_clk));
Sub0000000002  u_0000000066_Sub0000000002(.i_data_1(B[12][2]), .i_data_2(C[12][2]), .o_data(mult_result_i[12][2]), .i_clk(i_clk));
Sub0000000002  u_0000000067_Sub0000000002(.i_data_1(A[12][3]), .i_data_2(B[12][3]), .o_data(mult_result_r[12][3]), .i_clk(i_clk));
Sub0000000002  u_0000000068_Sub0000000002(.i_data_1(B[12][3]), .i_data_2(C[12][3]), .o_data(mult_result_i[12][3]), .i_clk(i_clk));
Sub0000000002  u_0000000069_Sub0000000002(.i_data_1(A[13][0]), .i_data_2(B[13][0]), .o_data(mult_result_r[13][0]), .i_clk(i_clk));
Sub0000000002  u_000000006A_Sub0000000002(.i_data_1(B[13][0]), .i_data_2(C[13][0]), .o_data(mult_result_i[13][0]), .i_clk(i_clk));
Sub0000000002  u_000000006B_Sub0000000002(.i_data_1(A[13][1]), .i_data_2(B[13][1]), .o_data(mult_result_r[13][1]), .i_clk(i_clk));
Sub0000000002  u_000000006C_Sub0000000002(.i_data_1(B[13][1]), .i_data_2(C[13][1]), .o_data(mult_result_i[13][1]), .i_clk(i_clk));
Sub0000000002  u_000000006D_Sub0000000002(.i_data_1(A[13][2]), .i_data_2(B[13][2]), .o_data(mult_result_r[13][2]), .i_clk(i_clk));
Sub0000000002  u_000000006E_Sub0000000002(.i_data_1(B[13][2]), .i_data_2(C[13][2]), .o_data(mult_result_i[13][2]), .i_clk(i_clk));
Sub0000000002  u_000000006F_Sub0000000002(.i_data_1(A[13][3]), .i_data_2(B[13][3]), .o_data(mult_result_r[13][3]), .i_clk(i_clk));
Sub0000000002  u_0000000070_Sub0000000002(.i_data_1(B[13][3]), .i_data_2(C[13][3]), .o_data(mult_result_i[13][3]), .i_clk(i_clk));
Sub0000000002  u_0000000071_Sub0000000002(.i_data_1(A[14][0]), .i_data_2(B[14][0]), .o_data(mult_result_r[14][0]), .i_clk(i_clk));
Sub0000000002  u_0000000072_Sub0000000002(.i_data_1(B[14][0]), .i_data_2(C[14][0]), .o_data(mult_result_i[14][0]), .i_clk(i_clk));
Sub0000000002  u_0000000073_Sub0000000002(.i_data_1(A[14][1]), .i_data_2(B[14][1]), .o_data(mult_result_r[14][1]), .i_clk(i_clk));
Sub0000000002  u_0000000074_Sub0000000002(.i_data_1(B[14][1]), .i_data_2(C[14][1]), .o_data(mult_result_i[14][1]), .i_clk(i_clk));
Sub0000000002  u_0000000075_Sub0000000002(.i_data_1(A[14][2]), .i_data_2(B[14][2]), .o_data(mult_result_r[14][2]), .i_clk(i_clk));
Sub0000000002  u_0000000076_Sub0000000002(.i_data_1(B[14][2]), .i_data_2(C[14][2]), .o_data(mult_result_i[14][2]), .i_clk(i_clk));
Sub0000000002  u_0000000077_Sub0000000002(.i_data_1(A[14][3]), .i_data_2(B[14][3]), .o_data(mult_result_r[14][3]), .i_clk(i_clk));
Sub0000000002  u_0000000078_Sub0000000002(.i_data_1(B[14][3]), .i_data_2(C[14][3]), .o_data(mult_result_i[14][3]), .i_clk(i_clk));
Sub0000000002  u_0000000079_Sub0000000002(.i_data_1(A[15][0]), .i_data_2(B[15][0]), .o_data(mult_result_r[15][0]), .i_clk(i_clk));
Sub0000000002  u_000000007A_Sub0000000002(.i_data_1(B[15][0]), .i_data_2(C[15][0]), .o_data(mult_result_i[15][0]), .i_clk(i_clk));
Sub0000000002  u_000000007B_Sub0000000002(.i_data_1(A[15][1]), .i_data_2(B[15][1]), .o_data(mult_result_r[15][1]), .i_clk(i_clk));
Sub0000000002  u_000000007C_Sub0000000002(.i_data_1(B[15][1]), .i_data_2(C[15][1]), .o_data(mult_result_i[15][1]), .i_clk(i_clk));
Sub0000000002  u_000000007D_Sub0000000002(.i_data_1(A[15][2]), .i_data_2(B[15][2]), .o_data(mult_result_r[15][2]), .i_clk(i_clk));
Sub0000000002  u_000000007E_Sub0000000002(.i_data_1(B[15][2]), .i_data_2(C[15][2]), .o_data(mult_result_i[15][2]), .i_clk(i_clk));
Sub0000000002  u_000000007F_Sub0000000002(.i_data_1(A[15][3]), .i_data_2(B[15][3]), .o_data(mult_result_r[15][3]), .i_clk(i_clk));
Sub0000000002  u_0000000080_Sub0000000002(.i_data_1(B[15][3]), .i_data_2(C[15][3]), .o_data(mult_result_i[15][3]), .i_clk(i_clk));
Sub0000000002  u_0000000081_Sub0000000002(.i_data_1(A[16][0]), .i_data_2(B[16][0]), .o_data(mult_result_r[16][0]), .i_clk(i_clk));
Sub0000000002  u_0000000082_Sub0000000002(.i_data_1(B[16][0]), .i_data_2(C[16][0]), .o_data(mult_result_i[16][0]), .i_clk(i_clk));
Sub0000000002  u_0000000083_Sub0000000002(.i_data_1(A[16][1]), .i_data_2(B[16][1]), .o_data(mult_result_r[16][1]), .i_clk(i_clk));
Sub0000000002  u_0000000084_Sub0000000002(.i_data_1(B[16][1]), .i_data_2(C[16][1]), .o_data(mult_result_i[16][1]), .i_clk(i_clk));
Sub0000000002  u_0000000085_Sub0000000002(.i_data_1(A[16][2]), .i_data_2(B[16][2]), .o_data(mult_result_r[16][2]), .i_clk(i_clk));
Sub0000000002  u_0000000086_Sub0000000002(.i_data_1(B[16][2]), .i_data_2(C[16][2]), .o_data(mult_result_i[16][2]), .i_clk(i_clk));
Sub0000000002  u_0000000087_Sub0000000002(.i_data_1(A[16][3]), .i_data_2(B[16][3]), .o_data(mult_result_r[16][3]), .i_clk(i_clk));
Sub0000000002  u_0000000088_Sub0000000002(.i_data_1(B[16][3]), .i_data_2(C[16][3]), .o_data(mult_result_i[16][3]), .i_clk(i_clk));
Sub0000000002  u_0000000089_Sub0000000002(.i_data_1(A[17][0]), .i_data_2(B[17][0]), .o_data(mult_result_r[17][0]), .i_clk(i_clk));
Sub0000000002  u_000000008A_Sub0000000002(.i_data_1(B[17][0]), .i_data_2(C[17][0]), .o_data(mult_result_i[17][0]), .i_clk(i_clk));
Sub0000000002  u_000000008B_Sub0000000002(.i_data_1(A[17][1]), .i_data_2(B[17][1]), .o_data(mult_result_r[17][1]), .i_clk(i_clk));
Sub0000000002  u_000000008C_Sub0000000002(.i_data_1(B[17][1]), .i_data_2(C[17][1]), .o_data(mult_result_i[17][1]), .i_clk(i_clk));
Sub0000000002  u_000000008D_Sub0000000002(.i_data_1(A[17][2]), .i_data_2(B[17][2]), .o_data(mult_result_r[17][2]), .i_clk(i_clk));
Sub0000000002  u_000000008E_Sub0000000002(.i_data_1(B[17][2]), .i_data_2(C[17][2]), .o_data(mult_result_i[17][2]), .i_clk(i_clk));
Sub0000000002  u_000000008F_Sub0000000002(.i_data_1(A[17][3]), .i_data_2(B[17][3]), .o_data(mult_result_r[17][3]), .i_clk(i_clk));
Sub0000000002  u_0000000090_Sub0000000002(.i_data_1(B[17][3]), .i_data_2(C[17][3]), .o_data(mult_result_i[17][3]), .i_clk(i_clk));
Sub0000000002  u_0000000091_Sub0000000002(.i_data_1(A[18][0]), .i_data_2(B[18][0]), .o_data(mult_result_r[18][0]), .i_clk(i_clk));
Sub0000000002  u_0000000092_Sub0000000002(.i_data_1(B[18][0]), .i_data_2(C[18][0]), .o_data(mult_result_i[18][0]), .i_clk(i_clk));
Sub0000000002  u_0000000093_Sub0000000002(.i_data_1(A[18][1]), .i_data_2(B[18][1]), .o_data(mult_result_r[18][1]), .i_clk(i_clk));
Sub0000000002  u_0000000094_Sub0000000002(.i_data_1(B[18][1]), .i_data_2(C[18][1]), .o_data(mult_result_i[18][1]), .i_clk(i_clk));
Sub0000000002  u_0000000095_Sub0000000002(.i_data_1(A[18][2]), .i_data_2(B[18][2]), .o_data(mult_result_r[18][2]), .i_clk(i_clk));
Sub0000000002  u_0000000096_Sub0000000002(.i_data_1(B[18][2]), .i_data_2(C[18][2]), .o_data(mult_result_i[18][2]), .i_clk(i_clk));
Sub0000000002  u_0000000097_Sub0000000002(.i_data_1(A[18][3]), .i_data_2(B[18][3]), .o_data(mult_result_r[18][3]), .i_clk(i_clk));
Sub0000000002  u_0000000098_Sub0000000002(.i_data_1(B[18][3]), .i_data_2(C[18][3]), .o_data(mult_result_i[18][3]), .i_clk(i_clk));
Sub0000000002  u_0000000099_Sub0000000002(.i_data_1(A[19][0]), .i_data_2(B[19][0]), .o_data(mult_result_r[19][0]), .i_clk(i_clk));
Sub0000000002  u_000000009A_Sub0000000002(.i_data_1(B[19][0]), .i_data_2(C[19][0]), .o_data(mult_result_i[19][0]), .i_clk(i_clk));
Sub0000000002  u_000000009B_Sub0000000002(.i_data_1(A[19][1]), .i_data_2(B[19][1]), .o_data(mult_result_r[19][1]), .i_clk(i_clk));
Sub0000000002  u_000000009C_Sub0000000002(.i_data_1(B[19][1]), .i_data_2(C[19][1]), .o_data(mult_result_i[19][1]), .i_clk(i_clk));
Sub0000000002  u_000000009D_Sub0000000002(.i_data_1(A[19][2]), .i_data_2(B[19][2]), .o_data(mult_result_r[19][2]), .i_clk(i_clk));
Sub0000000002  u_000000009E_Sub0000000002(.i_data_1(B[19][2]), .i_data_2(C[19][2]), .o_data(mult_result_i[19][2]), .i_clk(i_clk));
Sub0000000002  u_000000009F_Sub0000000002(.i_data_1(A[19][3]), .i_data_2(B[19][3]), .o_data(mult_result_r[19][3]), .i_clk(i_clk));
Sub0000000002  u_00000000A0_Sub0000000002(.i_data_1(B[19][3]), .i_data_2(C[19][3]), .o_data(mult_result_i[19][3]), .i_clk(i_clk));
Sub0000000002  u_00000000A1_Sub0000000002(.i_data_1(A[20][0]), .i_data_2(B[20][0]), .o_data(mult_result_r[20][0]), .i_clk(i_clk));
Sub0000000002  u_00000000A2_Sub0000000002(.i_data_1(B[20][0]), .i_data_2(C[20][0]), .o_data(mult_result_i[20][0]), .i_clk(i_clk));
Sub0000000002  u_00000000A3_Sub0000000002(.i_data_1(A[20][1]), .i_data_2(B[20][1]), .o_data(mult_result_r[20][1]), .i_clk(i_clk));
Sub0000000002  u_00000000A4_Sub0000000002(.i_data_1(B[20][1]), .i_data_2(C[20][1]), .o_data(mult_result_i[20][1]), .i_clk(i_clk));
Sub0000000002  u_00000000A5_Sub0000000002(.i_data_1(A[20][2]), .i_data_2(B[20][2]), .o_data(mult_result_r[20][2]), .i_clk(i_clk));
Sub0000000002  u_00000000A6_Sub0000000002(.i_data_1(B[20][2]), .i_data_2(C[20][2]), .o_data(mult_result_i[20][2]), .i_clk(i_clk));
Sub0000000002  u_00000000A7_Sub0000000002(.i_data_1(A[20][3]), .i_data_2(B[20][3]), .o_data(mult_result_r[20][3]), .i_clk(i_clk));
Sub0000000002  u_00000000A8_Sub0000000002(.i_data_1(B[20][3]), .i_data_2(C[20][3]), .o_data(mult_result_i[20][3]), .i_clk(i_clk));
Sub0000000002  u_00000000A9_Sub0000000002(.i_data_1(A[21][0]), .i_data_2(B[21][0]), .o_data(mult_result_r[21][0]), .i_clk(i_clk));
Sub0000000002  u_00000000AA_Sub0000000002(.i_data_1(B[21][0]), .i_data_2(C[21][0]), .o_data(mult_result_i[21][0]), .i_clk(i_clk));
Sub0000000002  u_00000000AB_Sub0000000002(.i_data_1(A[21][1]), .i_data_2(B[21][1]), .o_data(mult_result_r[21][1]), .i_clk(i_clk));
Sub0000000002  u_00000000AC_Sub0000000002(.i_data_1(B[21][1]), .i_data_2(C[21][1]), .o_data(mult_result_i[21][1]), .i_clk(i_clk));
Sub0000000002  u_00000000AD_Sub0000000002(.i_data_1(A[21][2]), .i_data_2(B[21][2]), .o_data(mult_result_r[21][2]), .i_clk(i_clk));
Sub0000000002  u_00000000AE_Sub0000000002(.i_data_1(B[21][2]), .i_data_2(C[21][2]), .o_data(mult_result_i[21][2]), .i_clk(i_clk));
Sub0000000002  u_00000000AF_Sub0000000002(.i_data_1(A[21][3]), .i_data_2(B[21][3]), .o_data(mult_result_r[21][3]), .i_clk(i_clk));
Sub0000000002  u_00000000B0_Sub0000000002(.i_data_1(B[21][3]), .i_data_2(C[21][3]), .o_data(mult_result_i[21][3]), .i_clk(i_clk));
Sub0000000002  u_00000000B1_Sub0000000002(.i_data_1(A[22][0]), .i_data_2(B[22][0]), .o_data(mult_result_r[22][0]), .i_clk(i_clk));
Sub0000000002  u_00000000B2_Sub0000000002(.i_data_1(B[22][0]), .i_data_2(C[22][0]), .o_data(mult_result_i[22][0]), .i_clk(i_clk));
Sub0000000002  u_00000000B3_Sub0000000002(.i_data_1(A[22][1]), .i_data_2(B[22][1]), .o_data(mult_result_r[22][1]), .i_clk(i_clk));
Sub0000000002  u_00000000B4_Sub0000000002(.i_data_1(B[22][1]), .i_data_2(C[22][1]), .o_data(mult_result_i[22][1]), .i_clk(i_clk));
Sub0000000002  u_00000000B5_Sub0000000002(.i_data_1(A[22][2]), .i_data_2(B[22][2]), .o_data(mult_result_r[22][2]), .i_clk(i_clk));
Sub0000000002  u_00000000B6_Sub0000000002(.i_data_1(B[22][2]), .i_data_2(C[22][2]), .o_data(mult_result_i[22][2]), .i_clk(i_clk));
Sub0000000002  u_00000000B7_Sub0000000002(.i_data_1(A[22][3]), .i_data_2(B[22][3]), .o_data(mult_result_r[22][3]), .i_clk(i_clk));
Sub0000000002  u_00000000B8_Sub0000000002(.i_data_1(B[22][3]), .i_data_2(C[22][3]), .o_data(mult_result_i[22][3]), .i_clk(i_clk));
Sub0000000002  u_00000000B9_Sub0000000002(.i_data_1(A[23][0]), .i_data_2(B[23][0]), .o_data(mult_result_r[23][0]), .i_clk(i_clk));
Sub0000000002  u_00000000BA_Sub0000000002(.i_data_1(B[23][0]), .i_data_2(C[23][0]), .o_data(mult_result_i[23][0]), .i_clk(i_clk));
Sub0000000002  u_00000000BB_Sub0000000002(.i_data_1(A[23][1]), .i_data_2(B[23][1]), .o_data(mult_result_r[23][1]), .i_clk(i_clk));
Sub0000000002  u_00000000BC_Sub0000000002(.i_data_1(B[23][1]), .i_data_2(C[23][1]), .o_data(mult_result_i[23][1]), .i_clk(i_clk));
Sub0000000002  u_00000000BD_Sub0000000002(.i_data_1(A[23][2]), .i_data_2(B[23][2]), .o_data(mult_result_r[23][2]), .i_clk(i_clk));
Sub0000000002  u_00000000BE_Sub0000000002(.i_data_1(B[23][2]), .i_data_2(C[23][2]), .o_data(mult_result_i[23][2]), .i_clk(i_clk));
Sub0000000002  u_00000000BF_Sub0000000002(.i_data_1(A[23][3]), .i_data_2(B[23][3]), .o_data(mult_result_r[23][3]), .i_clk(i_clk));
Sub0000000002  u_00000000C0_Sub0000000002(.i_data_1(B[23][3]), .i_data_2(C[23][3]), .o_data(mult_result_i[23][3]), .i_clk(i_clk));
Sub0000000002  u_00000000C1_Sub0000000002(.i_data_1(A[24][0]), .i_data_2(B[24][0]), .o_data(mult_result_r[24][0]), .i_clk(i_clk));
Sub0000000002  u_00000000C2_Sub0000000002(.i_data_1(B[24][0]), .i_data_2(C[24][0]), .o_data(mult_result_i[24][0]), .i_clk(i_clk));
Sub0000000002  u_00000000C3_Sub0000000002(.i_data_1(A[24][1]), .i_data_2(B[24][1]), .o_data(mult_result_r[24][1]), .i_clk(i_clk));
Sub0000000002  u_00000000C4_Sub0000000002(.i_data_1(B[24][1]), .i_data_2(C[24][1]), .o_data(mult_result_i[24][1]), .i_clk(i_clk));
Sub0000000002  u_00000000C5_Sub0000000002(.i_data_1(A[24][2]), .i_data_2(B[24][2]), .o_data(mult_result_r[24][2]), .i_clk(i_clk));
Sub0000000002  u_00000000C6_Sub0000000002(.i_data_1(B[24][2]), .i_data_2(C[24][2]), .o_data(mult_result_i[24][2]), .i_clk(i_clk));
Sub0000000002  u_00000000C7_Sub0000000002(.i_data_1(A[24][3]), .i_data_2(B[24][3]), .o_data(mult_result_r[24][3]), .i_clk(i_clk));
Sub0000000002  u_00000000C8_Sub0000000002(.i_data_1(B[24][3]), .i_data_2(C[24][3]), .o_data(mult_result_i[24][3]), .i_clk(i_clk));
Sub0000000002  u_00000000C9_Sub0000000002(.i_data_1(A[25][0]), .i_data_2(B[25][0]), .o_data(mult_result_r[25][0]), .i_clk(i_clk));
Sub0000000002  u_00000000CA_Sub0000000002(.i_data_1(B[25][0]), .i_data_2(C[25][0]), .o_data(mult_result_i[25][0]), .i_clk(i_clk));
Sub0000000002  u_00000000CB_Sub0000000002(.i_data_1(A[25][1]), .i_data_2(B[25][1]), .o_data(mult_result_r[25][1]), .i_clk(i_clk));
Sub0000000002  u_00000000CC_Sub0000000002(.i_data_1(B[25][1]), .i_data_2(C[25][1]), .o_data(mult_result_i[25][1]), .i_clk(i_clk));
Sub0000000002  u_00000000CD_Sub0000000002(.i_data_1(A[25][2]), .i_data_2(B[25][2]), .o_data(mult_result_r[25][2]), .i_clk(i_clk));
Sub0000000002  u_00000000CE_Sub0000000002(.i_data_1(B[25][2]), .i_data_2(C[25][2]), .o_data(mult_result_i[25][2]), .i_clk(i_clk));
Sub0000000002  u_00000000CF_Sub0000000002(.i_data_1(A[25][3]), .i_data_2(B[25][3]), .o_data(mult_result_r[25][3]), .i_clk(i_clk));
Sub0000000002  u_00000000D0_Sub0000000002(.i_data_1(B[25][3]), .i_data_2(C[25][3]), .o_data(mult_result_i[25][3]), .i_clk(i_clk));
Sub0000000002  u_00000000D1_Sub0000000002(.i_data_1(A[26][0]), .i_data_2(B[26][0]), .o_data(mult_result_r[26][0]), .i_clk(i_clk));
Sub0000000002  u_00000000D2_Sub0000000002(.i_data_1(B[26][0]), .i_data_2(C[26][0]), .o_data(mult_result_i[26][0]), .i_clk(i_clk));
Sub0000000002  u_00000000D3_Sub0000000002(.i_data_1(A[26][1]), .i_data_2(B[26][1]), .o_data(mult_result_r[26][1]), .i_clk(i_clk));
Sub0000000002  u_00000000D4_Sub0000000002(.i_data_1(B[26][1]), .i_data_2(C[26][1]), .o_data(mult_result_i[26][1]), .i_clk(i_clk));
Sub0000000002  u_00000000D5_Sub0000000002(.i_data_1(A[26][2]), .i_data_2(B[26][2]), .o_data(mult_result_r[26][2]), .i_clk(i_clk));
Sub0000000002  u_00000000D6_Sub0000000002(.i_data_1(B[26][2]), .i_data_2(C[26][2]), .o_data(mult_result_i[26][2]), .i_clk(i_clk));
Sub0000000002  u_00000000D7_Sub0000000002(.i_data_1(A[26][3]), .i_data_2(B[26][3]), .o_data(mult_result_r[26][3]), .i_clk(i_clk));
Sub0000000002  u_00000000D8_Sub0000000002(.i_data_1(B[26][3]), .i_data_2(C[26][3]), .o_data(mult_result_i[26][3]), .i_clk(i_clk));
Sub0000000002  u_00000000D9_Sub0000000002(.i_data_1(A[27][0]), .i_data_2(B[27][0]), .o_data(mult_result_r[27][0]), .i_clk(i_clk));
Sub0000000002  u_00000000DA_Sub0000000002(.i_data_1(B[27][0]), .i_data_2(C[27][0]), .o_data(mult_result_i[27][0]), .i_clk(i_clk));
Sub0000000002  u_00000000DB_Sub0000000002(.i_data_1(A[27][1]), .i_data_2(B[27][1]), .o_data(mult_result_r[27][1]), .i_clk(i_clk));
Sub0000000002  u_00000000DC_Sub0000000002(.i_data_1(B[27][1]), .i_data_2(C[27][1]), .o_data(mult_result_i[27][1]), .i_clk(i_clk));
Sub0000000002  u_00000000DD_Sub0000000002(.i_data_1(A[27][2]), .i_data_2(B[27][2]), .o_data(mult_result_r[27][2]), .i_clk(i_clk));
Sub0000000002  u_00000000DE_Sub0000000002(.i_data_1(B[27][2]), .i_data_2(C[27][2]), .o_data(mult_result_i[27][2]), .i_clk(i_clk));
Sub0000000002  u_00000000DF_Sub0000000002(.i_data_1(A[27][3]), .i_data_2(B[27][3]), .o_data(mult_result_r[27][3]), .i_clk(i_clk));
Sub0000000002  u_00000000E0_Sub0000000002(.i_data_1(B[27][3]), .i_data_2(C[27][3]), .o_data(mult_result_i[27][3]), .i_clk(i_clk));
Sub0000000002  u_00000000E1_Sub0000000002(.i_data_1(A[28][0]), .i_data_2(B[28][0]), .o_data(mult_result_r[28][0]), .i_clk(i_clk));
Sub0000000002  u_00000000E2_Sub0000000002(.i_data_1(B[28][0]), .i_data_2(C[28][0]), .o_data(mult_result_i[28][0]), .i_clk(i_clk));
Sub0000000002  u_00000000E3_Sub0000000002(.i_data_1(A[28][1]), .i_data_2(B[28][1]), .o_data(mult_result_r[28][1]), .i_clk(i_clk));
Sub0000000002  u_00000000E4_Sub0000000002(.i_data_1(B[28][1]), .i_data_2(C[28][1]), .o_data(mult_result_i[28][1]), .i_clk(i_clk));
Sub0000000002  u_00000000E5_Sub0000000002(.i_data_1(A[28][2]), .i_data_2(B[28][2]), .o_data(mult_result_r[28][2]), .i_clk(i_clk));
Sub0000000002  u_00000000E6_Sub0000000002(.i_data_1(B[28][2]), .i_data_2(C[28][2]), .o_data(mult_result_i[28][2]), .i_clk(i_clk));
Sub0000000002  u_00000000E7_Sub0000000002(.i_data_1(A[28][3]), .i_data_2(B[28][3]), .o_data(mult_result_r[28][3]), .i_clk(i_clk));
Sub0000000002  u_00000000E8_Sub0000000002(.i_data_1(B[28][3]), .i_data_2(C[28][3]), .o_data(mult_result_i[28][3]), .i_clk(i_clk));
Sub0000000002  u_00000000E9_Sub0000000002(.i_data_1(A[29][0]), .i_data_2(B[29][0]), .o_data(mult_result_r[29][0]), .i_clk(i_clk));
Sub0000000002  u_00000000EA_Sub0000000002(.i_data_1(B[29][0]), .i_data_2(C[29][0]), .o_data(mult_result_i[29][0]), .i_clk(i_clk));
Sub0000000002  u_00000000EB_Sub0000000002(.i_data_1(A[29][1]), .i_data_2(B[29][1]), .o_data(mult_result_r[29][1]), .i_clk(i_clk));
Sub0000000002  u_00000000EC_Sub0000000002(.i_data_1(B[29][1]), .i_data_2(C[29][1]), .o_data(mult_result_i[29][1]), .i_clk(i_clk));
Sub0000000002  u_00000000ED_Sub0000000002(.i_data_1(A[29][2]), .i_data_2(B[29][2]), .o_data(mult_result_r[29][2]), .i_clk(i_clk));
Sub0000000002  u_00000000EE_Sub0000000002(.i_data_1(B[29][2]), .i_data_2(C[29][2]), .o_data(mult_result_i[29][2]), .i_clk(i_clk));
Sub0000000002  u_00000000EF_Sub0000000002(.i_data_1(A[29][3]), .i_data_2(B[29][3]), .o_data(mult_result_r[29][3]), .i_clk(i_clk));
Sub0000000002  u_00000000F0_Sub0000000002(.i_data_1(B[29][3]), .i_data_2(C[29][3]), .o_data(mult_result_i[29][3]), .i_clk(i_clk));
Sub0000000002  u_00000000F1_Sub0000000002(.i_data_1(A[30][0]), .i_data_2(B[30][0]), .o_data(mult_result_r[30][0]), .i_clk(i_clk));
Sub0000000002  u_00000000F2_Sub0000000002(.i_data_1(B[30][0]), .i_data_2(C[30][0]), .o_data(mult_result_i[30][0]), .i_clk(i_clk));
Sub0000000002  u_00000000F3_Sub0000000002(.i_data_1(A[30][1]), .i_data_2(B[30][1]), .o_data(mult_result_r[30][1]), .i_clk(i_clk));
Sub0000000002  u_00000000F4_Sub0000000002(.i_data_1(B[30][1]), .i_data_2(C[30][1]), .o_data(mult_result_i[30][1]), .i_clk(i_clk));
Sub0000000002  u_00000000F5_Sub0000000002(.i_data_1(A[30][2]), .i_data_2(B[30][2]), .o_data(mult_result_r[30][2]), .i_clk(i_clk));
Sub0000000002  u_00000000F6_Sub0000000002(.i_data_1(B[30][2]), .i_data_2(C[30][2]), .o_data(mult_result_i[30][2]), .i_clk(i_clk));
Sub0000000002  u_00000000F7_Sub0000000002(.i_data_1(A[30][3]), .i_data_2(B[30][3]), .o_data(mult_result_r[30][3]), .i_clk(i_clk));
Sub0000000002  u_00000000F8_Sub0000000002(.i_data_1(B[30][3]), .i_data_2(C[30][3]), .o_data(mult_result_i[30][3]), .i_clk(i_clk));
Sub0000000002  u_00000000F9_Sub0000000002(.i_data_1(A[31][0]), .i_data_2(B[31][0]), .o_data(mult_result_r[31][0]), .i_clk(i_clk));
Sub0000000002  u_00000000FA_Sub0000000002(.i_data_1(B[31][0]), .i_data_2(C[31][0]), .o_data(mult_result_i[31][0]), .i_clk(i_clk));
Sub0000000002  u_00000000FB_Sub0000000002(.i_data_1(A[31][1]), .i_data_2(B[31][1]), .o_data(mult_result_r[31][1]), .i_clk(i_clk));
Sub0000000002  u_00000000FC_Sub0000000002(.i_data_1(B[31][1]), .i_data_2(C[31][1]), .o_data(mult_result_i[31][1]), .i_clk(i_clk));
Sub0000000002  u_00000000FD_Sub0000000002(.i_data_1(A[31][2]), .i_data_2(B[31][2]), .o_data(mult_result_r[31][2]), .i_clk(i_clk));
Sub0000000002  u_00000000FE_Sub0000000002(.i_data_1(B[31][2]), .i_data_2(C[31][2]), .o_data(mult_result_i[31][2]), .i_clk(i_clk));
Sub0000000002  u_00000000FF_Sub0000000002(.i_data_1(A[31][3]), .i_data_2(B[31][3]), .o_data(mult_result_r[31][3]), .i_clk(i_clk));
Sub0000000002  u_0000000100_Sub0000000002(.i_data_1(B[31][3]), .i_data_2(C[31][3]), .o_data(mult_result_i[31][3]), .i_clk(i_clk));
Sub0000000002  u_0000000101_Sub0000000002(.i_data_1(A[32][0]), .i_data_2(B[32][0]), .o_data(mult_result_r[32][0]), .i_clk(i_clk));
Sub0000000002  u_0000000102_Sub0000000002(.i_data_1(B[32][0]), .i_data_2(C[32][0]), .o_data(mult_result_i[32][0]), .i_clk(i_clk));
Sub0000000002  u_0000000103_Sub0000000002(.i_data_1(A[32][1]), .i_data_2(B[32][1]), .o_data(mult_result_r[32][1]), .i_clk(i_clk));
Sub0000000002  u_0000000104_Sub0000000002(.i_data_1(B[32][1]), .i_data_2(C[32][1]), .o_data(mult_result_i[32][1]), .i_clk(i_clk));
Sub0000000002  u_0000000105_Sub0000000002(.i_data_1(A[32][2]), .i_data_2(B[32][2]), .o_data(mult_result_r[32][2]), .i_clk(i_clk));
Sub0000000002  u_0000000106_Sub0000000002(.i_data_1(B[32][2]), .i_data_2(C[32][2]), .o_data(mult_result_i[32][2]), .i_clk(i_clk));
Sub0000000002  u_0000000107_Sub0000000002(.i_data_1(A[32][3]), .i_data_2(B[32][3]), .o_data(mult_result_r[32][3]), .i_clk(i_clk));
Sub0000000002  u_0000000108_Sub0000000002(.i_data_1(B[32][3]), .i_data_2(C[32][3]), .o_data(mult_result_i[32][3]), .i_clk(i_clk));
Sub0000000002  u_0000000109_Sub0000000002(.i_data_1(A[33][0]), .i_data_2(B[33][0]), .o_data(mult_result_r[33][0]), .i_clk(i_clk));
Sub0000000002  u_000000010A_Sub0000000002(.i_data_1(B[33][0]), .i_data_2(C[33][0]), .o_data(mult_result_i[33][0]), .i_clk(i_clk));
Sub0000000002  u_000000010B_Sub0000000002(.i_data_1(A[33][1]), .i_data_2(B[33][1]), .o_data(mult_result_r[33][1]), .i_clk(i_clk));
Sub0000000002  u_000000010C_Sub0000000002(.i_data_1(B[33][1]), .i_data_2(C[33][1]), .o_data(mult_result_i[33][1]), .i_clk(i_clk));
Sub0000000002  u_000000010D_Sub0000000002(.i_data_1(A[33][2]), .i_data_2(B[33][2]), .o_data(mult_result_r[33][2]), .i_clk(i_clk));
Sub0000000002  u_000000010E_Sub0000000002(.i_data_1(B[33][2]), .i_data_2(C[33][2]), .o_data(mult_result_i[33][2]), .i_clk(i_clk));
Sub0000000002  u_000000010F_Sub0000000002(.i_data_1(A[33][3]), .i_data_2(B[33][3]), .o_data(mult_result_r[33][3]), .i_clk(i_clk));
Sub0000000002  u_0000000110_Sub0000000002(.i_data_1(B[33][3]), .i_data_2(C[33][3]), .o_data(mult_result_i[33][3]), .i_clk(i_clk));
Sub0000000002  u_0000000111_Sub0000000002(.i_data_1(A[34][0]), .i_data_2(B[34][0]), .o_data(mult_result_r[34][0]), .i_clk(i_clk));
Sub0000000002  u_0000000112_Sub0000000002(.i_data_1(B[34][0]), .i_data_2(C[34][0]), .o_data(mult_result_i[34][0]), .i_clk(i_clk));
Sub0000000002  u_0000000113_Sub0000000002(.i_data_1(A[34][1]), .i_data_2(B[34][1]), .o_data(mult_result_r[34][1]), .i_clk(i_clk));
Sub0000000002  u_0000000114_Sub0000000002(.i_data_1(B[34][1]), .i_data_2(C[34][1]), .o_data(mult_result_i[34][1]), .i_clk(i_clk));
Sub0000000002  u_0000000115_Sub0000000002(.i_data_1(A[34][2]), .i_data_2(B[34][2]), .o_data(mult_result_r[34][2]), .i_clk(i_clk));
Sub0000000002  u_0000000116_Sub0000000002(.i_data_1(B[34][2]), .i_data_2(C[34][2]), .o_data(mult_result_i[34][2]), .i_clk(i_clk));
Sub0000000002  u_0000000117_Sub0000000002(.i_data_1(A[34][3]), .i_data_2(B[34][3]), .o_data(mult_result_r[34][3]), .i_clk(i_clk));
Sub0000000002  u_0000000118_Sub0000000002(.i_data_1(B[34][3]), .i_data_2(C[34][3]), .o_data(mult_result_i[34][3]), .i_clk(i_clk));
Sub0000000002  u_0000000119_Sub0000000002(.i_data_1(A[35][0]), .i_data_2(B[35][0]), .o_data(mult_result_r[35][0]), .i_clk(i_clk));
Sub0000000002  u_000000011A_Sub0000000002(.i_data_1(B[35][0]), .i_data_2(C[35][0]), .o_data(mult_result_i[35][0]), .i_clk(i_clk));
Sub0000000002  u_000000011B_Sub0000000002(.i_data_1(A[35][1]), .i_data_2(B[35][1]), .o_data(mult_result_r[35][1]), .i_clk(i_clk));
Sub0000000002  u_000000011C_Sub0000000002(.i_data_1(B[35][1]), .i_data_2(C[35][1]), .o_data(mult_result_i[35][1]), .i_clk(i_clk));
Sub0000000002  u_000000011D_Sub0000000002(.i_data_1(A[35][2]), .i_data_2(B[35][2]), .o_data(mult_result_r[35][2]), .i_clk(i_clk));
Sub0000000002  u_000000011E_Sub0000000002(.i_data_1(B[35][2]), .i_data_2(C[35][2]), .o_data(mult_result_i[35][2]), .i_clk(i_clk));
Sub0000000002  u_000000011F_Sub0000000002(.i_data_1(A[35][3]), .i_data_2(B[35][3]), .o_data(mult_result_r[35][3]), .i_clk(i_clk));
Sub0000000002  u_0000000120_Sub0000000002(.i_data_1(B[35][3]), .i_data_2(C[35][3]), .o_data(mult_result_i[35][3]), .i_clk(i_clk));
Sub0000000002  u_0000000121_Sub0000000002(.i_data_1(A[36][0]), .i_data_2(B[36][0]), .o_data(mult_result_r[36][0]), .i_clk(i_clk));
Sub0000000002  u_0000000122_Sub0000000002(.i_data_1(B[36][0]), .i_data_2(C[36][0]), .o_data(mult_result_i[36][0]), .i_clk(i_clk));
Sub0000000002  u_0000000123_Sub0000000002(.i_data_1(A[36][1]), .i_data_2(B[36][1]), .o_data(mult_result_r[36][1]), .i_clk(i_clk));
Sub0000000002  u_0000000124_Sub0000000002(.i_data_1(B[36][1]), .i_data_2(C[36][1]), .o_data(mult_result_i[36][1]), .i_clk(i_clk));
Sub0000000002  u_0000000125_Sub0000000002(.i_data_1(A[36][2]), .i_data_2(B[36][2]), .o_data(mult_result_r[36][2]), .i_clk(i_clk));
Sub0000000002  u_0000000126_Sub0000000002(.i_data_1(B[36][2]), .i_data_2(C[36][2]), .o_data(mult_result_i[36][2]), .i_clk(i_clk));
Sub0000000002  u_0000000127_Sub0000000002(.i_data_1(A[36][3]), .i_data_2(B[36][3]), .o_data(mult_result_r[36][3]), .i_clk(i_clk));
Sub0000000002  u_0000000128_Sub0000000002(.i_data_1(B[36][3]), .i_data_2(C[36][3]), .o_data(mult_result_i[36][3]), .i_clk(i_clk));
Sub0000000002  u_0000000129_Sub0000000002(.i_data_1(A[37][0]), .i_data_2(B[37][0]), .o_data(mult_result_r[37][0]), .i_clk(i_clk));
Sub0000000002  u_000000012A_Sub0000000002(.i_data_1(B[37][0]), .i_data_2(C[37][0]), .o_data(mult_result_i[37][0]), .i_clk(i_clk));
Sub0000000002  u_000000012B_Sub0000000002(.i_data_1(A[37][1]), .i_data_2(B[37][1]), .o_data(mult_result_r[37][1]), .i_clk(i_clk));
Sub0000000002  u_000000012C_Sub0000000002(.i_data_1(B[37][1]), .i_data_2(C[37][1]), .o_data(mult_result_i[37][1]), .i_clk(i_clk));
Sub0000000002  u_000000012D_Sub0000000002(.i_data_1(A[37][2]), .i_data_2(B[37][2]), .o_data(mult_result_r[37][2]), .i_clk(i_clk));
Sub0000000002  u_000000012E_Sub0000000002(.i_data_1(B[37][2]), .i_data_2(C[37][2]), .o_data(mult_result_i[37][2]), .i_clk(i_clk));
Sub0000000002  u_000000012F_Sub0000000002(.i_data_1(A[37][3]), .i_data_2(B[37][3]), .o_data(mult_result_r[37][3]), .i_clk(i_clk));
Sub0000000002  u_0000000130_Sub0000000002(.i_data_1(B[37][3]), .i_data_2(C[37][3]), .o_data(mult_result_i[37][3]), .i_clk(i_clk));
Sub0000000002  u_0000000131_Sub0000000002(.i_data_1(A[38][0]), .i_data_2(B[38][0]), .o_data(mult_result_r[38][0]), .i_clk(i_clk));
Sub0000000002  u_0000000132_Sub0000000002(.i_data_1(B[38][0]), .i_data_2(C[38][0]), .o_data(mult_result_i[38][0]), .i_clk(i_clk));
Sub0000000002  u_0000000133_Sub0000000002(.i_data_1(A[38][1]), .i_data_2(B[38][1]), .o_data(mult_result_r[38][1]), .i_clk(i_clk));
Sub0000000002  u_0000000134_Sub0000000002(.i_data_1(B[38][1]), .i_data_2(C[38][1]), .o_data(mult_result_i[38][1]), .i_clk(i_clk));
Sub0000000002  u_0000000135_Sub0000000002(.i_data_1(A[38][2]), .i_data_2(B[38][2]), .o_data(mult_result_r[38][2]), .i_clk(i_clk));
Sub0000000002  u_0000000136_Sub0000000002(.i_data_1(B[38][2]), .i_data_2(C[38][2]), .o_data(mult_result_i[38][2]), .i_clk(i_clk));
Sub0000000002  u_0000000137_Sub0000000002(.i_data_1(A[38][3]), .i_data_2(B[38][3]), .o_data(mult_result_r[38][3]), .i_clk(i_clk));
Sub0000000002  u_0000000138_Sub0000000002(.i_data_1(B[38][3]), .i_data_2(C[38][3]), .o_data(mult_result_i[38][3]), .i_clk(i_clk));
Sub0000000002  u_0000000139_Sub0000000002(.i_data_1(A[39][0]), .i_data_2(B[39][0]), .o_data(mult_result_r[39][0]), .i_clk(i_clk));
Sub0000000002  u_000000013A_Sub0000000002(.i_data_1(B[39][0]), .i_data_2(C[39][0]), .o_data(mult_result_i[39][0]), .i_clk(i_clk));
Sub0000000002  u_000000013B_Sub0000000002(.i_data_1(A[39][1]), .i_data_2(B[39][1]), .o_data(mult_result_r[39][1]), .i_clk(i_clk));
Sub0000000002  u_000000013C_Sub0000000002(.i_data_1(B[39][1]), .i_data_2(C[39][1]), .o_data(mult_result_i[39][1]), .i_clk(i_clk));
Sub0000000002  u_000000013D_Sub0000000002(.i_data_1(A[39][2]), .i_data_2(B[39][2]), .o_data(mult_result_r[39][2]), .i_clk(i_clk));
Sub0000000002  u_000000013E_Sub0000000002(.i_data_1(B[39][2]), .i_data_2(C[39][2]), .o_data(mult_result_i[39][2]), .i_clk(i_clk));
Sub0000000002  u_000000013F_Sub0000000002(.i_data_1(A[39][3]), .i_data_2(B[39][3]), .o_data(mult_result_r[39][3]), .i_clk(i_clk));
Sub0000000002  u_0000000140_Sub0000000002(.i_data_1(B[39][3]), .i_data_2(C[39][3]), .o_data(mult_result_i[39][3]), .i_clk(i_clk));
Sub0000000002  u_0000000141_Sub0000000002(.i_data_1(A[40][0]), .i_data_2(B[40][0]), .o_data(mult_result_r[40][0]), .i_clk(i_clk));
Sub0000000002  u_0000000142_Sub0000000002(.i_data_1(B[40][0]), .i_data_2(C[40][0]), .o_data(mult_result_i[40][0]), .i_clk(i_clk));
Sub0000000002  u_0000000143_Sub0000000002(.i_data_1(A[40][1]), .i_data_2(B[40][1]), .o_data(mult_result_r[40][1]), .i_clk(i_clk));
Sub0000000002  u_0000000144_Sub0000000002(.i_data_1(B[40][1]), .i_data_2(C[40][1]), .o_data(mult_result_i[40][1]), .i_clk(i_clk));
Sub0000000002  u_0000000145_Sub0000000002(.i_data_1(A[40][2]), .i_data_2(B[40][2]), .o_data(mult_result_r[40][2]), .i_clk(i_clk));
Sub0000000002  u_0000000146_Sub0000000002(.i_data_1(B[40][2]), .i_data_2(C[40][2]), .o_data(mult_result_i[40][2]), .i_clk(i_clk));
Sub0000000002  u_0000000147_Sub0000000002(.i_data_1(A[40][3]), .i_data_2(B[40][3]), .o_data(mult_result_r[40][3]), .i_clk(i_clk));
Sub0000000002  u_0000000148_Sub0000000002(.i_data_1(B[40][3]), .i_data_2(C[40][3]), .o_data(mult_result_i[40][3]), .i_clk(i_clk));
Sub0000000002  u_0000000149_Sub0000000002(.i_data_1(A[41][0]), .i_data_2(B[41][0]), .o_data(mult_result_r[41][0]), .i_clk(i_clk));
Sub0000000002  u_000000014A_Sub0000000002(.i_data_1(B[41][0]), .i_data_2(C[41][0]), .o_data(mult_result_i[41][0]), .i_clk(i_clk));
Sub0000000002  u_000000014B_Sub0000000002(.i_data_1(A[41][1]), .i_data_2(B[41][1]), .o_data(mult_result_r[41][1]), .i_clk(i_clk));
Sub0000000002  u_000000014C_Sub0000000002(.i_data_1(B[41][1]), .i_data_2(C[41][1]), .o_data(mult_result_i[41][1]), .i_clk(i_clk));
Sub0000000002  u_000000014D_Sub0000000002(.i_data_1(A[41][2]), .i_data_2(B[41][2]), .o_data(mult_result_r[41][2]), .i_clk(i_clk));
Sub0000000002  u_000000014E_Sub0000000002(.i_data_1(B[41][2]), .i_data_2(C[41][2]), .o_data(mult_result_i[41][2]), .i_clk(i_clk));
Sub0000000002  u_000000014F_Sub0000000002(.i_data_1(A[41][3]), .i_data_2(B[41][3]), .o_data(mult_result_r[41][3]), .i_clk(i_clk));
Sub0000000002  u_0000000150_Sub0000000002(.i_data_1(B[41][3]), .i_data_2(C[41][3]), .o_data(mult_result_i[41][3]), .i_clk(i_clk));
Sub0000000002  u_0000000151_Sub0000000002(.i_data_1(A[42][0]), .i_data_2(B[42][0]), .o_data(mult_result_r[42][0]), .i_clk(i_clk));
Sub0000000002  u_0000000152_Sub0000000002(.i_data_1(B[42][0]), .i_data_2(C[42][0]), .o_data(mult_result_i[42][0]), .i_clk(i_clk));
Sub0000000002  u_0000000153_Sub0000000002(.i_data_1(A[42][1]), .i_data_2(B[42][1]), .o_data(mult_result_r[42][1]), .i_clk(i_clk));
Sub0000000002  u_0000000154_Sub0000000002(.i_data_1(B[42][1]), .i_data_2(C[42][1]), .o_data(mult_result_i[42][1]), .i_clk(i_clk));
Sub0000000002  u_0000000155_Sub0000000002(.i_data_1(A[42][2]), .i_data_2(B[42][2]), .o_data(mult_result_r[42][2]), .i_clk(i_clk));
Sub0000000002  u_0000000156_Sub0000000002(.i_data_1(B[42][2]), .i_data_2(C[42][2]), .o_data(mult_result_i[42][2]), .i_clk(i_clk));
Sub0000000002  u_0000000157_Sub0000000002(.i_data_1(A[42][3]), .i_data_2(B[42][3]), .o_data(mult_result_r[42][3]), .i_clk(i_clk));
Sub0000000002  u_0000000158_Sub0000000002(.i_data_1(B[42][3]), .i_data_2(C[42][3]), .o_data(mult_result_i[42][3]), .i_clk(i_clk));
Sub0000000002  u_0000000159_Sub0000000002(.i_data_1(A[43][0]), .i_data_2(B[43][0]), .o_data(mult_result_r[43][0]), .i_clk(i_clk));
Sub0000000002  u_000000015A_Sub0000000002(.i_data_1(B[43][0]), .i_data_2(C[43][0]), .o_data(mult_result_i[43][0]), .i_clk(i_clk));
Sub0000000002  u_000000015B_Sub0000000002(.i_data_1(A[43][1]), .i_data_2(B[43][1]), .o_data(mult_result_r[43][1]), .i_clk(i_clk));
Sub0000000002  u_000000015C_Sub0000000002(.i_data_1(B[43][1]), .i_data_2(C[43][1]), .o_data(mult_result_i[43][1]), .i_clk(i_clk));
Sub0000000002  u_000000015D_Sub0000000002(.i_data_1(A[43][2]), .i_data_2(B[43][2]), .o_data(mult_result_r[43][2]), .i_clk(i_clk));
Sub0000000002  u_000000015E_Sub0000000002(.i_data_1(B[43][2]), .i_data_2(C[43][2]), .o_data(mult_result_i[43][2]), .i_clk(i_clk));
Sub0000000002  u_000000015F_Sub0000000002(.i_data_1(A[43][3]), .i_data_2(B[43][3]), .o_data(mult_result_r[43][3]), .i_clk(i_clk));
Sub0000000002  u_0000000160_Sub0000000002(.i_data_1(B[43][3]), .i_data_2(C[43][3]), .o_data(mult_result_i[43][3]), .i_clk(i_clk));
Sub0000000002  u_0000000161_Sub0000000002(.i_data_1(A[44][0]), .i_data_2(B[44][0]), .o_data(mult_result_r[44][0]), .i_clk(i_clk));
Sub0000000002  u_0000000162_Sub0000000002(.i_data_1(B[44][0]), .i_data_2(C[44][0]), .o_data(mult_result_i[44][0]), .i_clk(i_clk));
Sub0000000002  u_0000000163_Sub0000000002(.i_data_1(A[44][1]), .i_data_2(B[44][1]), .o_data(mult_result_r[44][1]), .i_clk(i_clk));
Sub0000000002  u_0000000164_Sub0000000002(.i_data_1(B[44][1]), .i_data_2(C[44][1]), .o_data(mult_result_i[44][1]), .i_clk(i_clk));
Sub0000000002  u_0000000165_Sub0000000002(.i_data_1(A[44][2]), .i_data_2(B[44][2]), .o_data(mult_result_r[44][2]), .i_clk(i_clk));
Sub0000000002  u_0000000166_Sub0000000002(.i_data_1(B[44][2]), .i_data_2(C[44][2]), .o_data(mult_result_i[44][2]), .i_clk(i_clk));
Sub0000000002  u_0000000167_Sub0000000002(.i_data_1(A[44][3]), .i_data_2(B[44][3]), .o_data(mult_result_r[44][3]), .i_clk(i_clk));
Sub0000000002  u_0000000168_Sub0000000002(.i_data_1(B[44][3]), .i_data_2(C[44][3]), .o_data(mult_result_i[44][3]), .i_clk(i_clk));
Sub0000000002  u_0000000169_Sub0000000002(.i_data_1(A[45][0]), .i_data_2(B[45][0]), .o_data(mult_result_r[45][0]), .i_clk(i_clk));
Sub0000000002  u_000000016A_Sub0000000002(.i_data_1(B[45][0]), .i_data_2(C[45][0]), .o_data(mult_result_i[45][0]), .i_clk(i_clk));
Sub0000000002  u_000000016B_Sub0000000002(.i_data_1(A[45][1]), .i_data_2(B[45][1]), .o_data(mult_result_r[45][1]), .i_clk(i_clk));
Sub0000000002  u_000000016C_Sub0000000002(.i_data_1(B[45][1]), .i_data_2(C[45][1]), .o_data(mult_result_i[45][1]), .i_clk(i_clk));
Sub0000000002  u_000000016D_Sub0000000002(.i_data_1(A[45][2]), .i_data_2(B[45][2]), .o_data(mult_result_r[45][2]), .i_clk(i_clk));
Sub0000000002  u_000000016E_Sub0000000002(.i_data_1(B[45][2]), .i_data_2(C[45][2]), .o_data(mult_result_i[45][2]), .i_clk(i_clk));
Sub0000000002  u_000000016F_Sub0000000002(.i_data_1(A[45][3]), .i_data_2(B[45][3]), .o_data(mult_result_r[45][3]), .i_clk(i_clk));
Sub0000000002  u_0000000170_Sub0000000002(.i_data_1(B[45][3]), .i_data_2(C[45][3]), .o_data(mult_result_i[45][3]), .i_clk(i_clk));
Sub0000000002  u_0000000171_Sub0000000002(.i_data_1(A[46][0]), .i_data_2(B[46][0]), .o_data(mult_result_r[46][0]), .i_clk(i_clk));
Sub0000000002  u_0000000172_Sub0000000002(.i_data_1(B[46][0]), .i_data_2(C[46][0]), .o_data(mult_result_i[46][0]), .i_clk(i_clk));
Sub0000000002  u_0000000173_Sub0000000002(.i_data_1(A[46][1]), .i_data_2(B[46][1]), .o_data(mult_result_r[46][1]), .i_clk(i_clk));
Sub0000000002  u_0000000174_Sub0000000002(.i_data_1(B[46][1]), .i_data_2(C[46][1]), .o_data(mult_result_i[46][1]), .i_clk(i_clk));
Sub0000000002  u_0000000175_Sub0000000002(.i_data_1(A[46][2]), .i_data_2(B[46][2]), .o_data(mult_result_r[46][2]), .i_clk(i_clk));
Sub0000000002  u_0000000176_Sub0000000002(.i_data_1(B[46][2]), .i_data_2(C[46][2]), .o_data(mult_result_i[46][2]), .i_clk(i_clk));
Sub0000000002  u_0000000177_Sub0000000002(.i_data_1(A[46][3]), .i_data_2(B[46][3]), .o_data(mult_result_r[46][3]), .i_clk(i_clk));
Sub0000000002  u_0000000178_Sub0000000002(.i_data_1(B[46][3]), .i_data_2(C[46][3]), .o_data(mult_result_i[46][3]), .i_clk(i_clk));
Sub0000000002  u_0000000179_Sub0000000002(.i_data_1(A[47][0]), .i_data_2(B[47][0]), .o_data(mult_result_r[47][0]), .i_clk(i_clk));
Sub0000000002  u_000000017A_Sub0000000002(.i_data_1(B[47][0]), .i_data_2(C[47][0]), .o_data(mult_result_i[47][0]), .i_clk(i_clk));
Sub0000000002  u_000000017B_Sub0000000002(.i_data_1(A[47][1]), .i_data_2(B[47][1]), .o_data(mult_result_r[47][1]), .i_clk(i_clk));
Sub0000000002  u_000000017C_Sub0000000002(.i_data_1(B[47][1]), .i_data_2(C[47][1]), .o_data(mult_result_i[47][1]), .i_clk(i_clk));
Sub0000000002  u_000000017D_Sub0000000002(.i_data_1(A[47][2]), .i_data_2(B[47][2]), .o_data(mult_result_r[47][2]), .i_clk(i_clk));
Sub0000000002  u_000000017E_Sub0000000002(.i_data_1(B[47][2]), .i_data_2(C[47][2]), .o_data(mult_result_i[47][2]), .i_clk(i_clk));
Sub0000000002  u_000000017F_Sub0000000002(.i_data_1(A[47][3]), .i_data_2(B[47][3]), .o_data(mult_result_r[47][3]), .i_clk(i_clk));
Sub0000000002  u_0000000180_Sub0000000002(.i_data_1(B[47][3]), .i_data_2(C[47][3]), .o_data(mult_result_i[47][3]), .i_clk(i_clk));
Sub0000000002  u_0000000181_Sub0000000002(.i_data_1(A[48][0]), .i_data_2(B[48][0]), .o_data(mult_result_r[48][0]), .i_clk(i_clk));
Sub0000000002  u_0000000182_Sub0000000002(.i_data_1(B[48][0]), .i_data_2(C[48][0]), .o_data(mult_result_i[48][0]), .i_clk(i_clk));
Sub0000000002  u_0000000183_Sub0000000002(.i_data_1(A[48][1]), .i_data_2(B[48][1]), .o_data(mult_result_r[48][1]), .i_clk(i_clk));
Sub0000000002  u_0000000184_Sub0000000002(.i_data_1(B[48][1]), .i_data_2(C[48][1]), .o_data(mult_result_i[48][1]), .i_clk(i_clk));
Sub0000000002  u_0000000185_Sub0000000002(.i_data_1(A[48][2]), .i_data_2(B[48][2]), .o_data(mult_result_r[48][2]), .i_clk(i_clk));
Sub0000000002  u_0000000186_Sub0000000002(.i_data_1(B[48][2]), .i_data_2(C[48][2]), .o_data(mult_result_i[48][2]), .i_clk(i_clk));
Sub0000000002  u_0000000187_Sub0000000002(.i_data_1(A[48][3]), .i_data_2(B[48][3]), .o_data(mult_result_r[48][3]), .i_clk(i_clk));
Sub0000000002  u_0000000188_Sub0000000002(.i_data_1(B[48][3]), .i_data_2(C[48][3]), .o_data(mult_result_i[48][3]), .i_clk(i_clk));
Sub0000000002  u_0000000189_Sub0000000002(.i_data_1(A[49][0]), .i_data_2(B[49][0]), .o_data(mult_result_r[49][0]), .i_clk(i_clk));
Sub0000000002  u_000000018A_Sub0000000002(.i_data_1(B[49][0]), .i_data_2(C[49][0]), .o_data(mult_result_i[49][0]), .i_clk(i_clk));
Sub0000000002  u_000000018B_Sub0000000002(.i_data_1(A[49][1]), .i_data_2(B[49][1]), .o_data(mult_result_r[49][1]), .i_clk(i_clk));
Sub0000000002  u_000000018C_Sub0000000002(.i_data_1(B[49][1]), .i_data_2(C[49][1]), .o_data(mult_result_i[49][1]), .i_clk(i_clk));
Sub0000000002  u_000000018D_Sub0000000002(.i_data_1(A[49][2]), .i_data_2(B[49][2]), .o_data(mult_result_r[49][2]), .i_clk(i_clk));
Sub0000000002  u_000000018E_Sub0000000002(.i_data_1(B[49][2]), .i_data_2(C[49][2]), .o_data(mult_result_i[49][2]), .i_clk(i_clk));
Sub0000000002  u_000000018F_Sub0000000002(.i_data_1(A[49][3]), .i_data_2(B[49][3]), .o_data(mult_result_r[49][3]), .i_clk(i_clk));
Sub0000000002  u_0000000190_Sub0000000002(.i_data_1(B[49][3]), .i_data_2(C[49][3]), .o_data(mult_result_i[49][3]), .i_clk(i_clk));
Sub0000000002  u_0000000191_Sub0000000002(.i_data_1(A[50][0]), .i_data_2(B[50][0]), .o_data(mult_result_r[50][0]), .i_clk(i_clk));
Sub0000000002  u_0000000192_Sub0000000002(.i_data_1(B[50][0]), .i_data_2(C[50][0]), .o_data(mult_result_i[50][0]), .i_clk(i_clk));
Sub0000000002  u_0000000193_Sub0000000002(.i_data_1(A[50][1]), .i_data_2(B[50][1]), .o_data(mult_result_r[50][1]), .i_clk(i_clk));
Sub0000000002  u_0000000194_Sub0000000002(.i_data_1(B[50][1]), .i_data_2(C[50][1]), .o_data(mult_result_i[50][1]), .i_clk(i_clk));
Sub0000000002  u_0000000195_Sub0000000002(.i_data_1(A[50][2]), .i_data_2(B[50][2]), .o_data(mult_result_r[50][2]), .i_clk(i_clk));
Sub0000000002  u_0000000196_Sub0000000002(.i_data_1(B[50][2]), .i_data_2(C[50][2]), .o_data(mult_result_i[50][2]), .i_clk(i_clk));
Sub0000000002  u_0000000197_Sub0000000002(.i_data_1(A[50][3]), .i_data_2(B[50][3]), .o_data(mult_result_r[50][3]), .i_clk(i_clk));
Sub0000000002  u_0000000198_Sub0000000002(.i_data_1(B[50][3]), .i_data_2(C[50][3]), .o_data(mult_result_i[50][3]), .i_clk(i_clk));
Sub0000000002  u_0000000199_Sub0000000002(.i_data_1(A[51][0]), .i_data_2(B[51][0]), .o_data(mult_result_r[51][0]), .i_clk(i_clk));
Sub0000000002  u_000000019A_Sub0000000002(.i_data_1(B[51][0]), .i_data_2(C[51][0]), .o_data(mult_result_i[51][0]), .i_clk(i_clk));
Sub0000000002  u_000000019B_Sub0000000002(.i_data_1(A[51][1]), .i_data_2(B[51][1]), .o_data(mult_result_r[51][1]), .i_clk(i_clk));
Sub0000000002  u_000000019C_Sub0000000002(.i_data_1(B[51][1]), .i_data_2(C[51][1]), .o_data(mult_result_i[51][1]), .i_clk(i_clk));
Sub0000000002  u_000000019D_Sub0000000002(.i_data_1(A[51][2]), .i_data_2(B[51][2]), .o_data(mult_result_r[51][2]), .i_clk(i_clk));
Sub0000000002  u_000000019E_Sub0000000002(.i_data_1(B[51][2]), .i_data_2(C[51][2]), .o_data(mult_result_i[51][2]), .i_clk(i_clk));
Sub0000000002  u_000000019F_Sub0000000002(.i_data_1(A[51][3]), .i_data_2(B[51][3]), .o_data(mult_result_r[51][3]), .i_clk(i_clk));
Sub0000000002  u_00000001A0_Sub0000000002(.i_data_1(B[51][3]), .i_data_2(C[51][3]), .o_data(mult_result_i[51][3]), .i_clk(i_clk));
Sub0000000002  u_00000001A1_Sub0000000002(.i_data_1(A[52][0]), .i_data_2(B[52][0]), .o_data(mult_result_r[52][0]), .i_clk(i_clk));
Sub0000000002  u_00000001A2_Sub0000000002(.i_data_1(B[52][0]), .i_data_2(C[52][0]), .o_data(mult_result_i[52][0]), .i_clk(i_clk));
Sub0000000002  u_00000001A3_Sub0000000002(.i_data_1(A[52][1]), .i_data_2(B[52][1]), .o_data(mult_result_r[52][1]), .i_clk(i_clk));
Sub0000000002  u_00000001A4_Sub0000000002(.i_data_1(B[52][1]), .i_data_2(C[52][1]), .o_data(mult_result_i[52][1]), .i_clk(i_clk));
Sub0000000002  u_00000001A5_Sub0000000002(.i_data_1(A[52][2]), .i_data_2(B[52][2]), .o_data(mult_result_r[52][2]), .i_clk(i_clk));
Sub0000000002  u_00000001A6_Sub0000000002(.i_data_1(B[52][2]), .i_data_2(C[52][2]), .o_data(mult_result_i[52][2]), .i_clk(i_clk));
Sub0000000002  u_00000001A7_Sub0000000002(.i_data_1(A[52][3]), .i_data_2(B[52][3]), .o_data(mult_result_r[52][3]), .i_clk(i_clk));
Sub0000000002  u_00000001A8_Sub0000000002(.i_data_1(B[52][3]), .i_data_2(C[52][3]), .o_data(mult_result_i[52][3]), .i_clk(i_clk));
Sub0000000002  u_00000001A9_Sub0000000002(.i_data_1(A[53][0]), .i_data_2(B[53][0]), .o_data(mult_result_r[53][0]), .i_clk(i_clk));
Sub0000000002  u_00000001AA_Sub0000000002(.i_data_1(B[53][0]), .i_data_2(C[53][0]), .o_data(mult_result_i[53][0]), .i_clk(i_clk));
Sub0000000002  u_00000001AB_Sub0000000002(.i_data_1(A[53][1]), .i_data_2(B[53][1]), .o_data(mult_result_r[53][1]), .i_clk(i_clk));
Sub0000000002  u_00000001AC_Sub0000000002(.i_data_1(B[53][1]), .i_data_2(C[53][1]), .o_data(mult_result_i[53][1]), .i_clk(i_clk));
Sub0000000002  u_00000001AD_Sub0000000002(.i_data_1(A[53][2]), .i_data_2(B[53][2]), .o_data(mult_result_r[53][2]), .i_clk(i_clk));
Sub0000000002  u_00000001AE_Sub0000000002(.i_data_1(B[53][2]), .i_data_2(C[53][2]), .o_data(mult_result_i[53][2]), .i_clk(i_clk));
Sub0000000002  u_00000001AF_Sub0000000002(.i_data_1(A[53][3]), .i_data_2(B[53][3]), .o_data(mult_result_r[53][3]), .i_clk(i_clk));
Sub0000000002  u_00000001B0_Sub0000000002(.i_data_1(B[53][3]), .i_data_2(C[53][3]), .o_data(mult_result_i[53][3]), .i_clk(i_clk));
Sub0000000002  u_00000001B1_Sub0000000002(.i_data_1(A[54][0]), .i_data_2(B[54][0]), .o_data(mult_result_r[54][0]), .i_clk(i_clk));
Sub0000000002  u_00000001B2_Sub0000000002(.i_data_1(B[54][0]), .i_data_2(C[54][0]), .o_data(mult_result_i[54][0]), .i_clk(i_clk));
Sub0000000002  u_00000001B3_Sub0000000002(.i_data_1(A[54][1]), .i_data_2(B[54][1]), .o_data(mult_result_r[54][1]), .i_clk(i_clk));
Sub0000000002  u_00000001B4_Sub0000000002(.i_data_1(B[54][1]), .i_data_2(C[54][1]), .o_data(mult_result_i[54][1]), .i_clk(i_clk));
Sub0000000002  u_00000001B5_Sub0000000002(.i_data_1(A[54][2]), .i_data_2(B[54][2]), .o_data(mult_result_r[54][2]), .i_clk(i_clk));
Sub0000000002  u_00000001B6_Sub0000000002(.i_data_1(B[54][2]), .i_data_2(C[54][2]), .o_data(mult_result_i[54][2]), .i_clk(i_clk));
Sub0000000002  u_00000001B7_Sub0000000002(.i_data_1(A[54][3]), .i_data_2(B[54][3]), .o_data(mult_result_r[54][3]), .i_clk(i_clk));
Sub0000000002  u_00000001B8_Sub0000000002(.i_data_1(B[54][3]), .i_data_2(C[54][3]), .o_data(mult_result_i[54][3]), .i_clk(i_clk));
Sub0000000002  u_00000001B9_Sub0000000002(.i_data_1(A[55][0]), .i_data_2(B[55][0]), .o_data(mult_result_r[55][0]), .i_clk(i_clk));
Sub0000000002  u_00000001BA_Sub0000000002(.i_data_1(B[55][0]), .i_data_2(C[55][0]), .o_data(mult_result_i[55][0]), .i_clk(i_clk));
Sub0000000002  u_00000001BB_Sub0000000002(.i_data_1(A[55][1]), .i_data_2(B[55][1]), .o_data(mult_result_r[55][1]), .i_clk(i_clk));
Sub0000000002  u_00000001BC_Sub0000000002(.i_data_1(B[55][1]), .i_data_2(C[55][1]), .o_data(mult_result_i[55][1]), .i_clk(i_clk));
Sub0000000002  u_00000001BD_Sub0000000002(.i_data_1(A[55][2]), .i_data_2(B[55][2]), .o_data(mult_result_r[55][2]), .i_clk(i_clk));
Sub0000000002  u_00000001BE_Sub0000000002(.i_data_1(B[55][2]), .i_data_2(C[55][2]), .o_data(mult_result_i[55][2]), .i_clk(i_clk));
Sub0000000002  u_00000001BF_Sub0000000002(.i_data_1(A[55][3]), .i_data_2(B[55][3]), .o_data(mult_result_r[55][3]), .i_clk(i_clk));
Sub0000000002  u_00000001C0_Sub0000000002(.i_data_1(B[55][3]), .i_data_2(C[55][3]), .o_data(mult_result_i[55][3]), .i_clk(i_clk));
Sub0000000002  u_00000001C1_Sub0000000002(.i_data_1(A[56][0]), .i_data_2(B[56][0]), .o_data(mult_result_r[56][0]), .i_clk(i_clk));
Sub0000000002  u_00000001C2_Sub0000000002(.i_data_1(B[56][0]), .i_data_2(C[56][0]), .o_data(mult_result_i[56][0]), .i_clk(i_clk));
Sub0000000002  u_00000001C3_Sub0000000002(.i_data_1(A[56][1]), .i_data_2(B[56][1]), .o_data(mult_result_r[56][1]), .i_clk(i_clk));
Sub0000000002  u_00000001C4_Sub0000000002(.i_data_1(B[56][1]), .i_data_2(C[56][1]), .o_data(mult_result_i[56][1]), .i_clk(i_clk));
Sub0000000002  u_00000001C5_Sub0000000002(.i_data_1(A[56][2]), .i_data_2(B[56][2]), .o_data(mult_result_r[56][2]), .i_clk(i_clk));
Sub0000000002  u_00000001C6_Sub0000000002(.i_data_1(B[56][2]), .i_data_2(C[56][2]), .o_data(mult_result_i[56][2]), .i_clk(i_clk));
Sub0000000002  u_00000001C7_Sub0000000002(.i_data_1(A[56][3]), .i_data_2(B[56][3]), .o_data(mult_result_r[56][3]), .i_clk(i_clk));
Sub0000000002  u_00000001C8_Sub0000000002(.i_data_1(B[56][3]), .i_data_2(C[56][3]), .o_data(mult_result_i[56][3]), .i_clk(i_clk));
Sub0000000002  u_00000001C9_Sub0000000002(.i_data_1(A[57][0]), .i_data_2(B[57][0]), .o_data(mult_result_r[57][0]), .i_clk(i_clk));
Sub0000000002  u_00000001CA_Sub0000000002(.i_data_1(B[57][0]), .i_data_2(C[57][0]), .o_data(mult_result_i[57][0]), .i_clk(i_clk));
Sub0000000002  u_00000001CB_Sub0000000002(.i_data_1(A[57][1]), .i_data_2(B[57][1]), .o_data(mult_result_r[57][1]), .i_clk(i_clk));
Sub0000000002  u_00000001CC_Sub0000000002(.i_data_1(B[57][1]), .i_data_2(C[57][1]), .o_data(mult_result_i[57][1]), .i_clk(i_clk));
Sub0000000002  u_00000001CD_Sub0000000002(.i_data_1(A[57][2]), .i_data_2(B[57][2]), .o_data(mult_result_r[57][2]), .i_clk(i_clk));
Sub0000000002  u_00000001CE_Sub0000000002(.i_data_1(B[57][2]), .i_data_2(C[57][2]), .o_data(mult_result_i[57][2]), .i_clk(i_clk));
Sub0000000002  u_00000001CF_Sub0000000002(.i_data_1(A[57][3]), .i_data_2(B[57][3]), .o_data(mult_result_r[57][3]), .i_clk(i_clk));
Sub0000000002  u_00000001D0_Sub0000000002(.i_data_1(B[57][3]), .i_data_2(C[57][3]), .o_data(mult_result_i[57][3]), .i_clk(i_clk));
Sub0000000002  u_00000001D1_Sub0000000002(.i_data_1(A[58][0]), .i_data_2(B[58][0]), .o_data(mult_result_r[58][0]), .i_clk(i_clk));
Sub0000000002  u_00000001D2_Sub0000000002(.i_data_1(B[58][0]), .i_data_2(C[58][0]), .o_data(mult_result_i[58][0]), .i_clk(i_clk));
Sub0000000002  u_00000001D3_Sub0000000002(.i_data_1(A[58][1]), .i_data_2(B[58][1]), .o_data(mult_result_r[58][1]), .i_clk(i_clk));
Sub0000000002  u_00000001D4_Sub0000000002(.i_data_1(B[58][1]), .i_data_2(C[58][1]), .o_data(mult_result_i[58][1]), .i_clk(i_clk));
Sub0000000002  u_00000001D5_Sub0000000002(.i_data_1(A[58][2]), .i_data_2(B[58][2]), .o_data(mult_result_r[58][2]), .i_clk(i_clk));
Sub0000000002  u_00000001D6_Sub0000000002(.i_data_1(B[58][2]), .i_data_2(C[58][2]), .o_data(mult_result_i[58][2]), .i_clk(i_clk));
Sub0000000002  u_00000001D7_Sub0000000002(.i_data_1(A[58][3]), .i_data_2(B[58][3]), .o_data(mult_result_r[58][3]), .i_clk(i_clk));
Sub0000000002  u_00000001D8_Sub0000000002(.i_data_1(B[58][3]), .i_data_2(C[58][3]), .o_data(mult_result_i[58][3]), .i_clk(i_clk));
Sub0000000002  u_00000001D9_Sub0000000002(.i_data_1(A[59][0]), .i_data_2(B[59][0]), .o_data(mult_result_r[59][0]), .i_clk(i_clk));
Sub0000000002  u_00000001DA_Sub0000000002(.i_data_1(B[59][0]), .i_data_2(C[59][0]), .o_data(mult_result_i[59][0]), .i_clk(i_clk));
Sub0000000002  u_00000001DB_Sub0000000002(.i_data_1(A[59][1]), .i_data_2(B[59][1]), .o_data(mult_result_r[59][1]), .i_clk(i_clk));
Sub0000000002  u_00000001DC_Sub0000000002(.i_data_1(B[59][1]), .i_data_2(C[59][1]), .o_data(mult_result_i[59][1]), .i_clk(i_clk));
Sub0000000002  u_00000001DD_Sub0000000002(.i_data_1(A[59][2]), .i_data_2(B[59][2]), .o_data(mult_result_r[59][2]), .i_clk(i_clk));
Sub0000000002  u_00000001DE_Sub0000000002(.i_data_1(B[59][2]), .i_data_2(C[59][2]), .o_data(mult_result_i[59][2]), .i_clk(i_clk));
Sub0000000002  u_00000001DF_Sub0000000002(.i_data_1(A[59][3]), .i_data_2(B[59][3]), .o_data(mult_result_r[59][3]), .i_clk(i_clk));
Sub0000000002  u_00000001E0_Sub0000000002(.i_data_1(B[59][3]), .i_data_2(C[59][3]), .o_data(mult_result_i[59][3]), .i_clk(i_clk));
Sub0000000002  u_00000001E1_Sub0000000002(.i_data_1(A[60][0]), .i_data_2(B[60][0]), .o_data(mult_result_r[60][0]), .i_clk(i_clk));
Sub0000000002  u_00000001E2_Sub0000000002(.i_data_1(B[60][0]), .i_data_2(C[60][0]), .o_data(mult_result_i[60][0]), .i_clk(i_clk));
Sub0000000002  u_00000001E3_Sub0000000002(.i_data_1(A[60][1]), .i_data_2(B[60][1]), .o_data(mult_result_r[60][1]), .i_clk(i_clk));
Sub0000000002  u_00000001E4_Sub0000000002(.i_data_1(B[60][1]), .i_data_2(C[60][1]), .o_data(mult_result_i[60][1]), .i_clk(i_clk));
Sub0000000002  u_00000001E5_Sub0000000002(.i_data_1(A[60][2]), .i_data_2(B[60][2]), .o_data(mult_result_r[60][2]), .i_clk(i_clk));
Sub0000000002  u_00000001E6_Sub0000000002(.i_data_1(B[60][2]), .i_data_2(C[60][2]), .o_data(mult_result_i[60][2]), .i_clk(i_clk));
Sub0000000002  u_00000001E7_Sub0000000002(.i_data_1(A[60][3]), .i_data_2(B[60][3]), .o_data(mult_result_r[60][3]), .i_clk(i_clk));
Sub0000000002  u_00000001E8_Sub0000000002(.i_data_1(B[60][3]), .i_data_2(C[60][3]), .o_data(mult_result_i[60][3]), .i_clk(i_clk));
Sub0000000002  u_00000001E9_Sub0000000002(.i_data_1(A[61][0]), .i_data_2(B[61][0]), .o_data(mult_result_r[61][0]), .i_clk(i_clk));
Sub0000000002  u_00000001EA_Sub0000000002(.i_data_1(B[61][0]), .i_data_2(C[61][0]), .o_data(mult_result_i[61][0]), .i_clk(i_clk));
Sub0000000002  u_00000001EB_Sub0000000002(.i_data_1(A[61][1]), .i_data_2(B[61][1]), .o_data(mult_result_r[61][1]), .i_clk(i_clk));
Sub0000000002  u_00000001EC_Sub0000000002(.i_data_1(B[61][1]), .i_data_2(C[61][1]), .o_data(mult_result_i[61][1]), .i_clk(i_clk));
Sub0000000002  u_00000001ED_Sub0000000002(.i_data_1(A[61][2]), .i_data_2(B[61][2]), .o_data(mult_result_r[61][2]), .i_clk(i_clk));
Sub0000000002  u_00000001EE_Sub0000000002(.i_data_1(B[61][2]), .i_data_2(C[61][2]), .o_data(mult_result_i[61][2]), .i_clk(i_clk));
Sub0000000002  u_00000001EF_Sub0000000002(.i_data_1(A[61][3]), .i_data_2(B[61][3]), .o_data(mult_result_r[61][3]), .i_clk(i_clk));
Sub0000000002  u_00000001F0_Sub0000000002(.i_data_1(B[61][3]), .i_data_2(C[61][3]), .o_data(mult_result_i[61][3]), .i_clk(i_clk));
Sub0000000002  u_00000001F1_Sub0000000002(.i_data_1(A[62][0]), .i_data_2(B[62][0]), .o_data(mult_result_r[62][0]), .i_clk(i_clk));
Sub0000000002  u_00000001F2_Sub0000000002(.i_data_1(B[62][0]), .i_data_2(C[62][0]), .o_data(mult_result_i[62][0]), .i_clk(i_clk));
Sub0000000002  u_00000001F3_Sub0000000002(.i_data_1(A[62][1]), .i_data_2(B[62][1]), .o_data(mult_result_r[62][1]), .i_clk(i_clk));
Sub0000000002  u_00000001F4_Sub0000000002(.i_data_1(B[62][1]), .i_data_2(C[62][1]), .o_data(mult_result_i[62][1]), .i_clk(i_clk));
Sub0000000002  u_00000001F5_Sub0000000002(.i_data_1(A[62][2]), .i_data_2(B[62][2]), .o_data(mult_result_r[62][2]), .i_clk(i_clk));
Sub0000000002  u_00000001F6_Sub0000000002(.i_data_1(B[62][2]), .i_data_2(C[62][2]), .o_data(mult_result_i[62][2]), .i_clk(i_clk));
Sub0000000002  u_00000001F7_Sub0000000002(.i_data_1(A[62][3]), .i_data_2(B[62][3]), .o_data(mult_result_r[62][3]), .i_clk(i_clk));
Sub0000000002  u_00000001F8_Sub0000000002(.i_data_1(B[62][3]), .i_data_2(C[62][3]), .o_data(mult_result_i[62][3]), .i_clk(i_clk));
Sub0000000002  u_00000001F9_Sub0000000002(.i_data_1(A[63][0]), .i_data_2(B[63][0]), .o_data(mult_result_r[63][0]), .i_clk(i_clk));
Sub0000000002  u_00000001FA_Sub0000000002(.i_data_1(B[63][0]), .i_data_2(C[63][0]), .o_data(mult_result_i[63][0]), .i_clk(i_clk));
Sub0000000002  u_00000001FB_Sub0000000002(.i_data_1(A[63][1]), .i_data_2(B[63][1]), .o_data(mult_result_r[63][1]), .i_clk(i_clk));
Sub0000000002  u_00000001FC_Sub0000000002(.i_data_1(B[63][1]), .i_data_2(C[63][1]), .o_data(mult_result_i[63][1]), .i_clk(i_clk));
Sub0000000002  u_00000001FD_Sub0000000002(.i_data_1(A[63][2]), .i_data_2(B[63][2]), .o_data(mult_result_r[63][2]), .i_clk(i_clk));
Sub0000000002  u_00000001FE_Sub0000000002(.i_data_1(B[63][2]), .i_data_2(C[63][2]), .o_data(mult_result_i[63][2]), .i_clk(i_clk));
Sub0000000002  u_00000001FF_Sub0000000002(.i_data_1(A[63][3]), .i_data_2(B[63][3]), .o_data(mult_result_r[63][3]), .i_clk(i_clk));
Sub0000000002  u_0000000200_Sub0000000002(.i_data_1(B[63][3]), .i_data_2(C[63][3]), .o_data(mult_result_i[63][3]), .i_clk(i_clk));
Sub0000000002  u_0000000201_Sub0000000002(.i_data_1(A[64][0]), .i_data_2(B[64][0]), .o_data(mult_result_r[64][0]), .i_clk(i_clk));
Sub0000000002  u_0000000202_Sub0000000002(.i_data_1(B[64][0]), .i_data_2(C[64][0]), .o_data(mult_result_i[64][0]), .i_clk(i_clk));
Sub0000000002  u_0000000203_Sub0000000002(.i_data_1(A[64][1]), .i_data_2(B[64][1]), .o_data(mult_result_r[64][1]), .i_clk(i_clk));
Sub0000000002  u_0000000204_Sub0000000002(.i_data_1(B[64][1]), .i_data_2(C[64][1]), .o_data(mult_result_i[64][1]), .i_clk(i_clk));
Sub0000000002  u_0000000205_Sub0000000002(.i_data_1(A[64][2]), .i_data_2(B[64][2]), .o_data(mult_result_r[64][2]), .i_clk(i_clk));
Sub0000000002  u_0000000206_Sub0000000002(.i_data_1(B[64][2]), .i_data_2(C[64][2]), .o_data(mult_result_i[64][2]), .i_clk(i_clk));
Sub0000000002  u_0000000207_Sub0000000002(.i_data_1(A[64][3]), .i_data_2(B[64][3]), .o_data(mult_result_r[64][3]), .i_clk(i_clk));
Sub0000000002  u_0000000208_Sub0000000002(.i_data_1(B[64][3]), .i_data_2(C[64][3]), .o_data(mult_result_i[64][3]), .i_clk(i_clk));
Sub0000000002  u_0000000209_Sub0000000002(.i_data_1(A[65][0]), .i_data_2(B[65][0]), .o_data(mult_result_r[65][0]), .i_clk(i_clk));
Sub0000000002  u_000000020A_Sub0000000002(.i_data_1(B[65][0]), .i_data_2(C[65][0]), .o_data(mult_result_i[65][0]), .i_clk(i_clk));
Sub0000000002  u_000000020B_Sub0000000002(.i_data_1(A[65][1]), .i_data_2(B[65][1]), .o_data(mult_result_r[65][1]), .i_clk(i_clk));
Sub0000000002  u_000000020C_Sub0000000002(.i_data_1(B[65][1]), .i_data_2(C[65][1]), .o_data(mult_result_i[65][1]), .i_clk(i_clk));
Sub0000000002  u_000000020D_Sub0000000002(.i_data_1(A[65][2]), .i_data_2(B[65][2]), .o_data(mult_result_r[65][2]), .i_clk(i_clk));
Sub0000000002  u_000000020E_Sub0000000002(.i_data_1(B[65][2]), .i_data_2(C[65][2]), .o_data(mult_result_i[65][2]), .i_clk(i_clk));
Sub0000000002  u_000000020F_Sub0000000002(.i_data_1(A[65][3]), .i_data_2(B[65][3]), .o_data(mult_result_r[65][3]), .i_clk(i_clk));
Sub0000000002  u_0000000210_Sub0000000002(.i_data_1(B[65][3]), .i_data_2(C[65][3]), .o_data(mult_result_i[65][3]), .i_clk(i_clk));
Sub0000000002  u_0000000211_Sub0000000002(.i_data_1(A[66][0]), .i_data_2(B[66][0]), .o_data(mult_result_r[66][0]), .i_clk(i_clk));
Sub0000000002  u_0000000212_Sub0000000002(.i_data_1(B[66][0]), .i_data_2(C[66][0]), .o_data(mult_result_i[66][0]), .i_clk(i_clk));
Sub0000000002  u_0000000213_Sub0000000002(.i_data_1(A[66][1]), .i_data_2(B[66][1]), .o_data(mult_result_r[66][1]), .i_clk(i_clk));
Sub0000000002  u_0000000214_Sub0000000002(.i_data_1(B[66][1]), .i_data_2(C[66][1]), .o_data(mult_result_i[66][1]), .i_clk(i_clk));
Sub0000000002  u_0000000215_Sub0000000002(.i_data_1(A[66][2]), .i_data_2(B[66][2]), .o_data(mult_result_r[66][2]), .i_clk(i_clk));
Sub0000000002  u_0000000216_Sub0000000002(.i_data_1(B[66][2]), .i_data_2(C[66][2]), .o_data(mult_result_i[66][2]), .i_clk(i_clk));
Sub0000000002  u_0000000217_Sub0000000002(.i_data_1(A[66][3]), .i_data_2(B[66][3]), .o_data(mult_result_r[66][3]), .i_clk(i_clk));
Sub0000000002  u_0000000218_Sub0000000002(.i_data_1(B[66][3]), .i_data_2(C[66][3]), .o_data(mult_result_i[66][3]), .i_clk(i_clk));
Sub0000000002  u_0000000219_Sub0000000002(.i_data_1(A[67][0]), .i_data_2(B[67][0]), .o_data(mult_result_r[67][0]), .i_clk(i_clk));
Sub0000000002  u_000000021A_Sub0000000002(.i_data_1(B[67][0]), .i_data_2(C[67][0]), .o_data(mult_result_i[67][0]), .i_clk(i_clk));
Sub0000000002  u_000000021B_Sub0000000002(.i_data_1(A[67][1]), .i_data_2(B[67][1]), .o_data(mult_result_r[67][1]), .i_clk(i_clk));
Sub0000000002  u_000000021C_Sub0000000002(.i_data_1(B[67][1]), .i_data_2(C[67][1]), .o_data(mult_result_i[67][1]), .i_clk(i_clk));
Sub0000000002  u_000000021D_Sub0000000002(.i_data_1(A[67][2]), .i_data_2(B[67][2]), .o_data(mult_result_r[67][2]), .i_clk(i_clk));
Sub0000000002  u_000000021E_Sub0000000002(.i_data_1(B[67][2]), .i_data_2(C[67][2]), .o_data(mult_result_i[67][2]), .i_clk(i_clk));
Sub0000000002  u_000000021F_Sub0000000002(.i_data_1(A[67][3]), .i_data_2(B[67][3]), .o_data(mult_result_r[67][3]), .i_clk(i_clk));
Sub0000000002  u_0000000220_Sub0000000002(.i_data_1(B[67][3]), .i_data_2(C[67][3]), .o_data(mult_result_i[67][3]), .i_clk(i_clk));
Sub0000000002  u_0000000221_Sub0000000002(.i_data_1(A[68][0]), .i_data_2(B[68][0]), .o_data(mult_result_r[68][0]), .i_clk(i_clk));
Sub0000000002  u_0000000222_Sub0000000002(.i_data_1(B[68][0]), .i_data_2(C[68][0]), .o_data(mult_result_i[68][0]), .i_clk(i_clk));
Sub0000000002  u_0000000223_Sub0000000002(.i_data_1(A[68][1]), .i_data_2(B[68][1]), .o_data(mult_result_r[68][1]), .i_clk(i_clk));
Sub0000000002  u_0000000224_Sub0000000002(.i_data_1(B[68][1]), .i_data_2(C[68][1]), .o_data(mult_result_i[68][1]), .i_clk(i_clk));
Sub0000000002  u_0000000225_Sub0000000002(.i_data_1(A[68][2]), .i_data_2(B[68][2]), .o_data(mult_result_r[68][2]), .i_clk(i_clk));
Sub0000000002  u_0000000226_Sub0000000002(.i_data_1(B[68][2]), .i_data_2(C[68][2]), .o_data(mult_result_i[68][2]), .i_clk(i_clk));
Sub0000000002  u_0000000227_Sub0000000002(.i_data_1(A[68][3]), .i_data_2(B[68][3]), .o_data(mult_result_r[68][3]), .i_clk(i_clk));
Sub0000000002  u_0000000228_Sub0000000002(.i_data_1(B[68][3]), .i_data_2(C[68][3]), .o_data(mult_result_i[68][3]), .i_clk(i_clk));
Sub0000000002  u_0000000229_Sub0000000002(.i_data_1(A[69][0]), .i_data_2(B[69][0]), .o_data(mult_result_r[69][0]), .i_clk(i_clk));
Sub0000000002  u_000000022A_Sub0000000002(.i_data_1(B[69][0]), .i_data_2(C[69][0]), .o_data(mult_result_i[69][0]), .i_clk(i_clk));
Sub0000000002  u_000000022B_Sub0000000002(.i_data_1(A[69][1]), .i_data_2(B[69][1]), .o_data(mult_result_r[69][1]), .i_clk(i_clk));
Sub0000000002  u_000000022C_Sub0000000002(.i_data_1(B[69][1]), .i_data_2(C[69][1]), .o_data(mult_result_i[69][1]), .i_clk(i_clk));
Sub0000000002  u_000000022D_Sub0000000002(.i_data_1(A[69][2]), .i_data_2(B[69][2]), .o_data(mult_result_r[69][2]), .i_clk(i_clk));
Sub0000000002  u_000000022E_Sub0000000002(.i_data_1(B[69][2]), .i_data_2(C[69][2]), .o_data(mult_result_i[69][2]), .i_clk(i_clk));
Sub0000000002  u_000000022F_Sub0000000002(.i_data_1(A[69][3]), .i_data_2(B[69][3]), .o_data(mult_result_r[69][3]), .i_clk(i_clk));
Sub0000000002  u_0000000230_Sub0000000002(.i_data_1(B[69][3]), .i_data_2(C[69][3]), .o_data(mult_result_i[69][3]), .i_clk(i_clk));
Sub0000000002  u_0000000231_Sub0000000002(.i_data_1(A[70][0]), .i_data_2(B[70][0]), .o_data(mult_result_r[70][0]), .i_clk(i_clk));
Sub0000000002  u_0000000232_Sub0000000002(.i_data_1(B[70][0]), .i_data_2(C[70][0]), .o_data(mult_result_i[70][0]), .i_clk(i_clk));
Sub0000000002  u_0000000233_Sub0000000002(.i_data_1(A[70][1]), .i_data_2(B[70][1]), .o_data(mult_result_r[70][1]), .i_clk(i_clk));
Sub0000000002  u_0000000234_Sub0000000002(.i_data_1(B[70][1]), .i_data_2(C[70][1]), .o_data(mult_result_i[70][1]), .i_clk(i_clk));
Sub0000000002  u_0000000235_Sub0000000002(.i_data_1(A[70][2]), .i_data_2(B[70][2]), .o_data(mult_result_r[70][2]), .i_clk(i_clk));
Sub0000000002  u_0000000236_Sub0000000002(.i_data_1(B[70][2]), .i_data_2(C[70][2]), .o_data(mult_result_i[70][2]), .i_clk(i_clk));
Sub0000000002  u_0000000237_Sub0000000002(.i_data_1(A[70][3]), .i_data_2(B[70][3]), .o_data(mult_result_r[70][3]), .i_clk(i_clk));
Sub0000000002  u_0000000238_Sub0000000002(.i_data_1(B[70][3]), .i_data_2(C[70][3]), .o_data(mult_result_i[70][3]), .i_clk(i_clk));
Sub0000000002  u_0000000239_Sub0000000002(.i_data_1(A[71][0]), .i_data_2(B[71][0]), .o_data(mult_result_r[71][0]), .i_clk(i_clk));
Sub0000000002  u_000000023A_Sub0000000002(.i_data_1(B[71][0]), .i_data_2(C[71][0]), .o_data(mult_result_i[71][0]), .i_clk(i_clk));
Sub0000000002  u_000000023B_Sub0000000002(.i_data_1(A[71][1]), .i_data_2(B[71][1]), .o_data(mult_result_r[71][1]), .i_clk(i_clk));
Sub0000000002  u_000000023C_Sub0000000002(.i_data_1(B[71][1]), .i_data_2(C[71][1]), .o_data(mult_result_i[71][1]), .i_clk(i_clk));
Sub0000000002  u_000000023D_Sub0000000002(.i_data_1(A[71][2]), .i_data_2(B[71][2]), .o_data(mult_result_r[71][2]), .i_clk(i_clk));
Sub0000000002  u_000000023E_Sub0000000002(.i_data_1(B[71][2]), .i_data_2(C[71][2]), .o_data(mult_result_i[71][2]), .i_clk(i_clk));
Sub0000000002  u_000000023F_Sub0000000002(.i_data_1(A[71][3]), .i_data_2(B[71][3]), .o_data(mult_result_r[71][3]), .i_clk(i_clk));
Sub0000000002  u_0000000240_Sub0000000002(.i_data_1(B[71][3]), .i_data_2(C[71][3]), .o_data(mult_result_i[71][3]), .i_clk(i_clk));
Sub0000000002  u_0000000241_Sub0000000002(.i_data_1(A[72][0]), .i_data_2(B[72][0]), .o_data(mult_result_r[72][0]), .i_clk(i_clk));
Sub0000000002  u_0000000242_Sub0000000002(.i_data_1(B[72][0]), .i_data_2(C[72][0]), .o_data(mult_result_i[72][0]), .i_clk(i_clk));
Sub0000000002  u_0000000243_Sub0000000002(.i_data_1(A[72][1]), .i_data_2(B[72][1]), .o_data(mult_result_r[72][1]), .i_clk(i_clk));
Sub0000000002  u_0000000244_Sub0000000002(.i_data_1(B[72][1]), .i_data_2(C[72][1]), .o_data(mult_result_i[72][1]), .i_clk(i_clk));
Sub0000000002  u_0000000245_Sub0000000002(.i_data_1(A[72][2]), .i_data_2(B[72][2]), .o_data(mult_result_r[72][2]), .i_clk(i_clk));
Sub0000000002  u_0000000246_Sub0000000002(.i_data_1(B[72][2]), .i_data_2(C[72][2]), .o_data(mult_result_i[72][2]), .i_clk(i_clk));
Sub0000000002  u_0000000247_Sub0000000002(.i_data_1(A[72][3]), .i_data_2(B[72][3]), .o_data(mult_result_r[72][3]), .i_clk(i_clk));
Sub0000000002  u_0000000248_Sub0000000002(.i_data_1(B[72][3]), .i_data_2(C[72][3]), .o_data(mult_result_i[72][3]), .i_clk(i_clk));
Sub0000000002  u_0000000249_Sub0000000002(.i_data_1(A[73][0]), .i_data_2(B[73][0]), .o_data(mult_result_r[73][0]), .i_clk(i_clk));
Sub0000000002  u_000000024A_Sub0000000002(.i_data_1(B[73][0]), .i_data_2(C[73][0]), .o_data(mult_result_i[73][0]), .i_clk(i_clk));
Sub0000000002  u_000000024B_Sub0000000002(.i_data_1(A[73][1]), .i_data_2(B[73][1]), .o_data(mult_result_r[73][1]), .i_clk(i_clk));
Sub0000000002  u_000000024C_Sub0000000002(.i_data_1(B[73][1]), .i_data_2(C[73][1]), .o_data(mult_result_i[73][1]), .i_clk(i_clk));
Sub0000000002  u_000000024D_Sub0000000002(.i_data_1(A[73][2]), .i_data_2(B[73][2]), .o_data(mult_result_r[73][2]), .i_clk(i_clk));
Sub0000000002  u_000000024E_Sub0000000002(.i_data_1(B[73][2]), .i_data_2(C[73][2]), .o_data(mult_result_i[73][2]), .i_clk(i_clk));
Sub0000000002  u_000000024F_Sub0000000002(.i_data_1(A[73][3]), .i_data_2(B[73][3]), .o_data(mult_result_r[73][3]), .i_clk(i_clk));
Sub0000000002  u_0000000250_Sub0000000002(.i_data_1(B[73][3]), .i_data_2(C[73][3]), .o_data(mult_result_i[73][3]), .i_clk(i_clk));
Sub0000000002  u_0000000251_Sub0000000002(.i_data_1(A[74][0]), .i_data_2(B[74][0]), .o_data(mult_result_r[74][0]), .i_clk(i_clk));
Sub0000000002  u_0000000252_Sub0000000002(.i_data_1(B[74][0]), .i_data_2(C[74][0]), .o_data(mult_result_i[74][0]), .i_clk(i_clk));
Sub0000000002  u_0000000253_Sub0000000002(.i_data_1(A[74][1]), .i_data_2(B[74][1]), .o_data(mult_result_r[74][1]), .i_clk(i_clk));
Sub0000000002  u_0000000254_Sub0000000002(.i_data_1(B[74][1]), .i_data_2(C[74][1]), .o_data(mult_result_i[74][1]), .i_clk(i_clk));
Sub0000000002  u_0000000255_Sub0000000002(.i_data_1(A[74][2]), .i_data_2(B[74][2]), .o_data(mult_result_r[74][2]), .i_clk(i_clk));
Sub0000000002  u_0000000256_Sub0000000002(.i_data_1(B[74][2]), .i_data_2(C[74][2]), .o_data(mult_result_i[74][2]), .i_clk(i_clk));
Sub0000000002  u_0000000257_Sub0000000002(.i_data_1(A[74][3]), .i_data_2(B[74][3]), .o_data(mult_result_r[74][3]), .i_clk(i_clk));
Sub0000000002  u_0000000258_Sub0000000002(.i_data_1(B[74][3]), .i_data_2(C[74][3]), .o_data(mult_result_i[74][3]), .i_clk(i_clk));
Sub0000000002  u_0000000259_Sub0000000002(.i_data_1(A[75][0]), .i_data_2(B[75][0]), .o_data(mult_result_r[75][0]), .i_clk(i_clk));
Sub0000000002  u_000000025A_Sub0000000002(.i_data_1(B[75][0]), .i_data_2(C[75][0]), .o_data(mult_result_i[75][0]), .i_clk(i_clk));
Sub0000000002  u_000000025B_Sub0000000002(.i_data_1(A[75][1]), .i_data_2(B[75][1]), .o_data(mult_result_r[75][1]), .i_clk(i_clk));
Sub0000000002  u_000000025C_Sub0000000002(.i_data_1(B[75][1]), .i_data_2(C[75][1]), .o_data(mult_result_i[75][1]), .i_clk(i_clk));
Sub0000000002  u_000000025D_Sub0000000002(.i_data_1(A[75][2]), .i_data_2(B[75][2]), .o_data(mult_result_r[75][2]), .i_clk(i_clk));
Sub0000000002  u_000000025E_Sub0000000002(.i_data_1(B[75][2]), .i_data_2(C[75][2]), .o_data(mult_result_i[75][2]), .i_clk(i_clk));
Sub0000000002  u_000000025F_Sub0000000002(.i_data_1(A[75][3]), .i_data_2(B[75][3]), .o_data(mult_result_r[75][3]), .i_clk(i_clk));
Sub0000000002  u_0000000260_Sub0000000002(.i_data_1(B[75][3]), .i_data_2(C[75][3]), .o_data(mult_result_i[75][3]), .i_clk(i_clk));
Sub0000000002  u_0000000261_Sub0000000002(.i_data_1(A[76][0]), .i_data_2(B[76][0]), .o_data(mult_result_r[76][0]), .i_clk(i_clk));
Sub0000000002  u_0000000262_Sub0000000002(.i_data_1(B[76][0]), .i_data_2(C[76][0]), .o_data(mult_result_i[76][0]), .i_clk(i_clk));
Sub0000000002  u_0000000263_Sub0000000002(.i_data_1(A[76][1]), .i_data_2(B[76][1]), .o_data(mult_result_r[76][1]), .i_clk(i_clk));
Sub0000000002  u_0000000264_Sub0000000002(.i_data_1(B[76][1]), .i_data_2(C[76][1]), .o_data(mult_result_i[76][1]), .i_clk(i_clk));
Sub0000000002  u_0000000265_Sub0000000002(.i_data_1(A[76][2]), .i_data_2(B[76][2]), .o_data(mult_result_r[76][2]), .i_clk(i_clk));
Sub0000000002  u_0000000266_Sub0000000002(.i_data_1(B[76][2]), .i_data_2(C[76][2]), .o_data(mult_result_i[76][2]), .i_clk(i_clk));
Sub0000000002  u_0000000267_Sub0000000002(.i_data_1(A[76][3]), .i_data_2(B[76][3]), .o_data(mult_result_r[76][3]), .i_clk(i_clk));
Sub0000000002  u_0000000268_Sub0000000002(.i_data_1(B[76][3]), .i_data_2(C[76][3]), .o_data(mult_result_i[76][3]), .i_clk(i_clk));
Sub0000000002  u_0000000269_Sub0000000002(.i_data_1(A[77][0]), .i_data_2(B[77][0]), .o_data(mult_result_r[77][0]), .i_clk(i_clk));
Sub0000000002  u_000000026A_Sub0000000002(.i_data_1(B[77][0]), .i_data_2(C[77][0]), .o_data(mult_result_i[77][0]), .i_clk(i_clk));
Sub0000000002  u_000000026B_Sub0000000002(.i_data_1(A[77][1]), .i_data_2(B[77][1]), .o_data(mult_result_r[77][1]), .i_clk(i_clk));
Sub0000000002  u_000000026C_Sub0000000002(.i_data_1(B[77][1]), .i_data_2(C[77][1]), .o_data(mult_result_i[77][1]), .i_clk(i_clk));
Sub0000000002  u_000000026D_Sub0000000002(.i_data_1(A[77][2]), .i_data_2(B[77][2]), .o_data(mult_result_r[77][2]), .i_clk(i_clk));
Sub0000000002  u_000000026E_Sub0000000002(.i_data_1(B[77][2]), .i_data_2(C[77][2]), .o_data(mult_result_i[77][2]), .i_clk(i_clk));
Sub0000000002  u_000000026F_Sub0000000002(.i_data_1(A[77][3]), .i_data_2(B[77][3]), .o_data(mult_result_r[77][3]), .i_clk(i_clk));
Sub0000000002  u_0000000270_Sub0000000002(.i_data_1(B[77][3]), .i_data_2(C[77][3]), .o_data(mult_result_i[77][3]), .i_clk(i_clk));
Sub0000000002  u_0000000271_Sub0000000002(.i_data_1(A[78][0]), .i_data_2(B[78][0]), .o_data(mult_result_r[78][0]), .i_clk(i_clk));
Sub0000000002  u_0000000272_Sub0000000002(.i_data_1(B[78][0]), .i_data_2(C[78][0]), .o_data(mult_result_i[78][0]), .i_clk(i_clk));
Sub0000000002  u_0000000273_Sub0000000002(.i_data_1(A[78][1]), .i_data_2(B[78][1]), .o_data(mult_result_r[78][1]), .i_clk(i_clk));
Sub0000000002  u_0000000274_Sub0000000002(.i_data_1(B[78][1]), .i_data_2(C[78][1]), .o_data(mult_result_i[78][1]), .i_clk(i_clk));
Sub0000000002  u_0000000275_Sub0000000002(.i_data_1(A[78][2]), .i_data_2(B[78][2]), .o_data(mult_result_r[78][2]), .i_clk(i_clk));
Sub0000000002  u_0000000276_Sub0000000002(.i_data_1(B[78][2]), .i_data_2(C[78][2]), .o_data(mult_result_i[78][2]), .i_clk(i_clk));
Sub0000000002  u_0000000277_Sub0000000002(.i_data_1(A[78][3]), .i_data_2(B[78][3]), .o_data(mult_result_r[78][3]), .i_clk(i_clk));
Sub0000000002  u_0000000278_Sub0000000002(.i_data_1(B[78][3]), .i_data_2(C[78][3]), .o_data(mult_result_i[78][3]), .i_clk(i_clk));
Sub0000000002  u_0000000279_Sub0000000002(.i_data_1(A[79][0]), .i_data_2(B[79][0]), .o_data(mult_result_r[79][0]), .i_clk(i_clk));
Sub0000000002  u_000000027A_Sub0000000002(.i_data_1(B[79][0]), .i_data_2(C[79][0]), .o_data(mult_result_i[79][0]), .i_clk(i_clk));
Sub0000000002  u_000000027B_Sub0000000002(.i_data_1(A[79][1]), .i_data_2(B[79][1]), .o_data(mult_result_r[79][1]), .i_clk(i_clk));
Sub0000000002  u_000000027C_Sub0000000002(.i_data_1(B[79][1]), .i_data_2(C[79][1]), .o_data(mult_result_i[79][1]), .i_clk(i_clk));
Sub0000000002  u_000000027D_Sub0000000002(.i_data_1(A[79][2]), .i_data_2(B[79][2]), .o_data(mult_result_r[79][2]), .i_clk(i_clk));
Sub0000000002  u_000000027E_Sub0000000002(.i_data_1(B[79][2]), .i_data_2(C[79][2]), .o_data(mult_result_i[79][2]), .i_clk(i_clk));
Sub0000000002  u_000000027F_Sub0000000002(.i_data_1(A[79][3]), .i_data_2(B[79][3]), .o_data(mult_result_r[79][3]), .i_clk(i_clk));
Sub0000000002  u_0000000280_Sub0000000002(.i_data_1(B[79][3]), .i_data_2(C[79][3]), .o_data(mult_result_i[79][3]), .i_clk(i_clk));
Sub0000000002  u_0000000281_Sub0000000002(.i_data_1(A[80][0]), .i_data_2(B[80][0]), .o_data(mult_result_r[80][0]), .i_clk(i_clk));
Sub0000000002  u_0000000282_Sub0000000002(.i_data_1(B[80][0]), .i_data_2(C[80][0]), .o_data(mult_result_i[80][0]), .i_clk(i_clk));
Sub0000000002  u_0000000283_Sub0000000002(.i_data_1(A[80][1]), .i_data_2(B[80][1]), .o_data(mult_result_r[80][1]), .i_clk(i_clk));
Sub0000000002  u_0000000284_Sub0000000002(.i_data_1(B[80][1]), .i_data_2(C[80][1]), .o_data(mult_result_i[80][1]), .i_clk(i_clk));
Sub0000000002  u_0000000285_Sub0000000002(.i_data_1(A[80][2]), .i_data_2(B[80][2]), .o_data(mult_result_r[80][2]), .i_clk(i_clk));
Sub0000000002  u_0000000286_Sub0000000002(.i_data_1(B[80][2]), .i_data_2(C[80][2]), .o_data(mult_result_i[80][2]), .i_clk(i_clk));
Sub0000000002  u_0000000287_Sub0000000002(.i_data_1(A[80][3]), .i_data_2(B[80][3]), .o_data(mult_result_r[80][3]), .i_clk(i_clk));
Sub0000000002  u_0000000288_Sub0000000002(.i_data_1(B[80][3]), .i_data_2(C[80][3]), .o_data(mult_result_i[80][3]), .i_clk(i_clk));
Sub0000000002  u_0000000289_Sub0000000002(.i_data_1(A[81][0]), .i_data_2(B[81][0]), .o_data(mult_result_r[81][0]), .i_clk(i_clk));
Sub0000000002  u_000000028A_Sub0000000002(.i_data_1(B[81][0]), .i_data_2(C[81][0]), .o_data(mult_result_i[81][0]), .i_clk(i_clk));
Sub0000000002  u_000000028B_Sub0000000002(.i_data_1(A[81][1]), .i_data_2(B[81][1]), .o_data(mult_result_r[81][1]), .i_clk(i_clk));
Sub0000000002  u_000000028C_Sub0000000002(.i_data_1(B[81][1]), .i_data_2(C[81][1]), .o_data(mult_result_i[81][1]), .i_clk(i_clk));
Sub0000000002  u_000000028D_Sub0000000002(.i_data_1(A[81][2]), .i_data_2(B[81][2]), .o_data(mult_result_r[81][2]), .i_clk(i_clk));
Sub0000000002  u_000000028E_Sub0000000002(.i_data_1(B[81][2]), .i_data_2(C[81][2]), .o_data(mult_result_i[81][2]), .i_clk(i_clk));
Sub0000000002  u_000000028F_Sub0000000002(.i_data_1(A[81][3]), .i_data_2(B[81][3]), .o_data(mult_result_r[81][3]), .i_clk(i_clk));
Sub0000000002  u_0000000290_Sub0000000002(.i_data_1(B[81][3]), .i_data_2(C[81][3]), .o_data(mult_result_i[81][3]), .i_clk(i_clk));
Sub0000000002  u_0000000291_Sub0000000002(.i_data_1(A[82][0]), .i_data_2(B[82][0]), .o_data(mult_result_r[82][0]), .i_clk(i_clk));
Sub0000000002  u_0000000292_Sub0000000002(.i_data_1(B[82][0]), .i_data_2(C[82][0]), .o_data(mult_result_i[82][0]), .i_clk(i_clk));
Sub0000000002  u_0000000293_Sub0000000002(.i_data_1(A[82][1]), .i_data_2(B[82][1]), .o_data(mult_result_r[82][1]), .i_clk(i_clk));
Sub0000000002  u_0000000294_Sub0000000002(.i_data_1(B[82][1]), .i_data_2(C[82][1]), .o_data(mult_result_i[82][1]), .i_clk(i_clk));
Sub0000000002  u_0000000295_Sub0000000002(.i_data_1(A[82][2]), .i_data_2(B[82][2]), .o_data(mult_result_r[82][2]), .i_clk(i_clk));
Sub0000000002  u_0000000296_Sub0000000002(.i_data_1(B[82][2]), .i_data_2(C[82][2]), .o_data(mult_result_i[82][2]), .i_clk(i_clk));
Sub0000000002  u_0000000297_Sub0000000002(.i_data_1(A[82][3]), .i_data_2(B[82][3]), .o_data(mult_result_r[82][3]), .i_clk(i_clk));
Sub0000000002  u_0000000298_Sub0000000002(.i_data_1(B[82][3]), .i_data_2(C[82][3]), .o_data(mult_result_i[82][3]), .i_clk(i_clk));
Sub0000000002  u_0000000299_Sub0000000002(.i_data_1(A[83][0]), .i_data_2(B[83][0]), .o_data(mult_result_r[83][0]), .i_clk(i_clk));
Sub0000000002  u_000000029A_Sub0000000002(.i_data_1(B[83][0]), .i_data_2(C[83][0]), .o_data(mult_result_i[83][0]), .i_clk(i_clk));
Sub0000000002  u_000000029B_Sub0000000002(.i_data_1(A[83][1]), .i_data_2(B[83][1]), .o_data(mult_result_r[83][1]), .i_clk(i_clk));
Sub0000000002  u_000000029C_Sub0000000002(.i_data_1(B[83][1]), .i_data_2(C[83][1]), .o_data(mult_result_i[83][1]), .i_clk(i_clk));
Sub0000000002  u_000000029D_Sub0000000002(.i_data_1(A[83][2]), .i_data_2(B[83][2]), .o_data(mult_result_r[83][2]), .i_clk(i_clk));
Sub0000000002  u_000000029E_Sub0000000002(.i_data_1(B[83][2]), .i_data_2(C[83][2]), .o_data(mult_result_i[83][2]), .i_clk(i_clk));
Sub0000000002  u_000000029F_Sub0000000002(.i_data_1(A[83][3]), .i_data_2(B[83][3]), .o_data(mult_result_r[83][3]), .i_clk(i_clk));
Sub0000000002  u_00000002A0_Sub0000000002(.i_data_1(B[83][3]), .i_data_2(C[83][3]), .o_data(mult_result_i[83][3]), .i_clk(i_clk));
Sub0000000002  u_00000002A1_Sub0000000002(.i_data_1(A[84][0]), .i_data_2(B[84][0]), .o_data(mult_result_r[84][0]), .i_clk(i_clk));
Sub0000000002  u_00000002A2_Sub0000000002(.i_data_1(B[84][0]), .i_data_2(C[84][0]), .o_data(mult_result_i[84][0]), .i_clk(i_clk));
Sub0000000002  u_00000002A3_Sub0000000002(.i_data_1(A[84][1]), .i_data_2(B[84][1]), .o_data(mult_result_r[84][1]), .i_clk(i_clk));
Sub0000000002  u_00000002A4_Sub0000000002(.i_data_1(B[84][1]), .i_data_2(C[84][1]), .o_data(mult_result_i[84][1]), .i_clk(i_clk));
Sub0000000002  u_00000002A5_Sub0000000002(.i_data_1(A[84][2]), .i_data_2(B[84][2]), .o_data(mult_result_r[84][2]), .i_clk(i_clk));
Sub0000000002  u_00000002A6_Sub0000000002(.i_data_1(B[84][2]), .i_data_2(C[84][2]), .o_data(mult_result_i[84][2]), .i_clk(i_clk));
Sub0000000002  u_00000002A7_Sub0000000002(.i_data_1(A[84][3]), .i_data_2(B[84][3]), .o_data(mult_result_r[84][3]), .i_clk(i_clk));
Sub0000000002  u_00000002A8_Sub0000000002(.i_data_1(B[84][3]), .i_data_2(C[84][3]), .o_data(mult_result_i[84][3]), .i_clk(i_clk));
Sub0000000002  u_00000002A9_Sub0000000002(.i_data_1(A[85][0]), .i_data_2(B[85][0]), .o_data(mult_result_r[85][0]), .i_clk(i_clk));
Sub0000000002  u_00000002AA_Sub0000000002(.i_data_1(B[85][0]), .i_data_2(C[85][0]), .o_data(mult_result_i[85][0]), .i_clk(i_clk));
Sub0000000002  u_00000002AB_Sub0000000002(.i_data_1(A[85][1]), .i_data_2(B[85][1]), .o_data(mult_result_r[85][1]), .i_clk(i_clk));
Sub0000000002  u_00000002AC_Sub0000000002(.i_data_1(B[85][1]), .i_data_2(C[85][1]), .o_data(mult_result_i[85][1]), .i_clk(i_clk));
Sub0000000002  u_00000002AD_Sub0000000002(.i_data_1(A[85][2]), .i_data_2(B[85][2]), .o_data(mult_result_r[85][2]), .i_clk(i_clk));
Sub0000000002  u_00000002AE_Sub0000000002(.i_data_1(B[85][2]), .i_data_2(C[85][2]), .o_data(mult_result_i[85][2]), .i_clk(i_clk));
Sub0000000002  u_00000002AF_Sub0000000002(.i_data_1(A[85][3]), .i_data_2(B[85][3]), .o_data(mult_result_r[85][3]), .i_clk(i_clk));
Sub0000000002  u_00000002B0_Sub0000000002(.i_data_1(B[85][3]), .i_data_2(C[85][3]), .o_data(mult_result_i[85][3]), .i_clk(i_clk));
Sub0000000002  u_00000002B1_Sub0000000002(.i_data_1(A[86][0]), .i_data_2(B[86][0]), .o_data(mult_result_r[86][0]), .i_clk(i_clk));
Sub0000000002  u_00000002B2_Sub0000000002(.i_data_1(B[86][0]), .i_data_2(C[86][0]), .o_data(mult_result_i[86][0]), .i_clk(i_clk));
Sub0000000002  u_00000002B3_Sub0000000002(.i_data_1(A[86][1]), .i_data_2(B[86][1]), .o_data(mult_result_r[86][1]), .i_clk(i_clk));
Sub0000000002  u_00000002B4_Sub0000000002(.i_data_1(B[86][1]), .i_data_2(C[86][1]), .o_data(mult_result_i[86][1]), .i_clk(i_clk));
Sub0000000002  u_00000002B5_Sub0000000002(.i_data_1(A[86][2]), .i_data_2(B[86][2]), .o_data(mult_result_r[86][2]), .i_clk(i_clk));
Sub0000000002  u_00000002B6_Sub0000000002(.i_data_1(B[86][2]), .i_data_2(C[86][2]), .o_data(mult_result_i[86][2]), .i_clk(i_clk));
Sub0000000002  u_00000002B7_Sub0000000002(.i_data_1(A[86][3]), .i_data_2(B[86][3]), .o_data(mult_result_r[86][3]), .i_clk(i_clk));
Sub0000000002  u_00000002B8_Sub0000000002(.i_data_1(B[86][3]), .i_data_2(C[86][3]), .o_data(mult_result_i[86][3]), .i_clk(i_clk));
Sub0000000002  u_00000002B9_Sub0000000002(.i_data_1(A[87][0]), .i_data_2(B[87][0]), .o_data(mult_result_r[87][0]), .i_clk(i_clk));
Sub0000000002  u_00000002BA_Sub0000000002(.i_data_1(B[87][0]), .i_data_2(C[87][0]), .o_data(mult_result_i[87][0]), .i_clk(i_clk));
Sub0000000002  u_00000002BB_Sub0000000002(.i_data_1(A[87][1]), .i_data_2(B[87][1]), .o_data(mult_result_r[87][1]), .i_clk(i_clk));
Sub0000000002  u_00000002BC_Sub0000000002(.i_data_1(B[87][1]), .i_data_2(C[87][1]), .o_data(mult_result_i[87][1]), .i_clk(i_clk));
Sub0000000002  u_00000002BD_Sub0000000002(.i_data_1(A[87][2]), .i_data_2(B[87][2]), .o_data(mult_result_r[87][2]), .i_clk(i_clk));
Sub0000000002  u_00000002BE_Sub0000000002(.i_data_1(B[87][2]), .i_data_2(C[87][2]), .o_data(mult_result_i[87][2]), .i_clk(i_clk));
Sub0000000002  u_00000002BF_Sub0000000002(.i_data_1(A[87][3]), .i_data_2(B[87][3]), .o_data(mult_result_r[87][3]), .i_clk(i_clk));
Sub0000000002  u_00000002C0_Sub0000000002(.i_data_1(B[87][3]), .i_data_2(C[87][3]), .o_data(mult_result_i[87][3]), .i_clk(i_clk));
Sub0000000002  u_00000002C1_Sub0000000002(.i_data_1(A[88][0]), .i_data_2(B[88][0]), .o_data(mult_result_r[88][0]), .i_clk(i_clk));
Sub0000000002  u_00000002C2_Sub0000000002(.i_data_1(B[88][0]), .i_data_2(C[88][0]), .o_data(mult_result_i[88][0]), .i_clk(i_clk));
Sub0000000002  u_00000002C3_Sub0000000002(.i_data_1(A[88][1]), .i_data_2(B[88][1]), .o_data(mult_result_r[88][1]), .i_clk(i_clk));
Sub0000000002  u_00000002C4_Sub0000000002(.i_data_1(B[88][1]), .i_data_2(C[88][1]), .o_data(mult_result_i[88][1]), .i_clk(i_clk));
Sub0000000002  u_00000002C5_Sub0000000002(.i_data_1(A[88][2]), .i_data_2(B[88][2]), .o_data(mult_result_r[88][2]), .i_clk(i_clk));
Sub0000000002  u_00000002C6_Sub0000000002(.i_data_1(B[88][2]), .i_data_2(C[88][2]), .o_data(mult_result_i[88][2]), .i_clk(i_clk));
Sub0000000002  u_00000002C7_Sub0000000002(.i_data_1(A[88][3]), .i_data_2(B[88][3]), .o_data(mult_result_r[88][3]), .i_clk(i_clk));
Sub0000000002  u_00000002C8_Sub0000000002(.i_data_1(B[88][3]), .i_data_2(C[88][3]), .o_data(mult_result_i[88][3]), .i_clk(i_clk));
Sub0000000002  u_00000002C9_Sub0000000002(.i_data_1(A[89][0]), .i_data_2(B[89][0]), .o_data(mult_result_r[89][0]), .i_clk(i_clk));
Sub0000000002  u_00000002CA_Sub0000000002(.i_data_1(B[89][0]), .i_data_2(C[89][0]), .o_data(mult_result_i[89][0]), .i_clk(i_clk));
Sub0000000002  u_00000002CB_Sub0000000002(.i_data_1(A[89][1]), .i_data_2(B[89][1]), .o_data(mult_result_r[89][1]), .i_clk(i_clk));
Sub0000000002  u_00000002CC_Sub0000000002(.i_data_1(B[89][1]), .i_data_2(C[89][1]), .o_data(mult_result_i[89][1]), .i_clk(i_clk));
Sub0000000002  u_00000002CD_Sub0000000002(.i_data_1(A[89][2]), .i_data_2(B[89][2]), .o_data(mult_result_r[89][2]), .i_clk(i_clk));
Sub0000000002  u_00000002CE_Sub0000000002(.i_data_1(B[89][2]), .i_data_2(C[89][2]), .o_data(mult_result_i[89][2]), .i_clk(i_clk));
Sub0000000002  u_00000002CF_Sub0000000002(.i_data_1(A[89][3]), .i_data_2(B[89][3]), .o_data(mult_result_r[89][3]), .i_clk(i_clk));
Sub0000000002  u_00000002D0_Sub0000000002(.i_data_1(B[89][3]), .i_data_2(C[89][3]), .o_data(mult_result_i[89][3]), .i_clk(i_clk));
Sub0000000002  u_00000002D1_Sub0000000002(.i_data_1(A[90][0]), .i_data_2(B[90][0]), .o_data(mult_result_r[90][0]), .i_clk(i_clk));
Sub0000000002  u_00000002D2_Sub0000000002(.i_data_1(B[90][0]), .i_data_2(C[90][0]), .o_data(mult_result_i[90][0]), .i_clk(i_clk));
Sub0000000002  u_00000002D3_Sub0000000002(.i_data_1(A[90][1]), .i_data_2(B[90][1]), .o_data(mult_result_r[90][1]), .i_clk(i_clk));
Sub0000000002  u_00000002D4_Sub0000000002(.i_data_1(B[90][1]), .i_data_2(C[90][1]), .o_data(mult_result_i[90][1]), .i_clk(i_clk));
Sub0000000002  u_00000002D5_Sub0000000002(.i_data_1(A[90][2]), .i_data_2(B[90][2]), .o_data(mult_result_r[90][2]), .i_clk(i_clk));
Sub0000000002  u_00000002D6_Sub0000000002(.i_data_1(B[90][2]), .i_data_2(C[90][2]), .o_data(mult_result_i[90][2]), .i_clk(i_clk));
Sub0000000002  u_00000002D7_Sub0000000002(.i_data_1(A[90][3]), .i_data_2(B[90][3]), .o_data(mult_result_r[90][3]), .i_clk(i_clk));
Sub0000000002  u_00000002D8_Sub0000000002(.i_data_1(B[90][3]), .i_data_2(C[90][3]), .o_data(mult_result_i[90][3]), .i_clk(i_clk));
Sub0000000002  u_00000002D9_Sub0000000002(.i_data_1(A[91][0]), .i_data_2(B[91][0]), .o_data(mult_result_r[91][0]), .i_clk(i_clk));
Sub0000000002  u_00000002DA_Sub0000000002(.i_data_1(B[91][0]), .i_data_2(C[91][0]), .o_data(mult_result_i[91][0]), .i_clk(i_clk));
Sub0000000002  u_00000002DB_Sub0000000002(.i_data_1(A[91][1]), .i_data_2(B[91][1]), .o_data(mult_result_r[91][1]), .i_clk(i_clk));
Sub0000000002  u_00000002DC_Sub0000000002(.i_data_1(B[91][1]), .i_data_2(C[91][1]), .o_data(mult_result_i[91][1]), .i_clk(i_clk));
Sub0000000002  u_00000002DD_Sub0000000002(.i_data_1(A[91][2]), .i_data_2(B[91][2]), .o_data(mult_result_r[91][2]), .i_clk(i_clk));
Sub0000000002  u_00000002DE_Sub0000000002(.i_data_1(B[91][2]), .i_data_2(C[91][2]), .o_data(mult_result_i[91][2]), .i_clk(i_clk));
Sub0000000002  u_00000002DF_Sub0000000002(.i_data_1(A[91][3]), .i_data_2(B[91][3]), .o_data(mult_result_r[91][3]), .i_clk(i_clk));
Sub0000000002  u_00000002E0_Sub0000000002(.i_data_1(B[91][3]), .i_data_2(C[91][3]), .o_data(mult_result_i[91][3]), .i_clk(i_clk));
Sub0000000002  u_00000002E1_Sub0000000002(.i_data_1(A[92][0]), .i_data_2(B[92][0]), .o_data(mult_result_r[92][0]), .i_clk(i_clk));
Sub0000000002  u_00000002E2_Sub0000000002(.i_data_1(B[92][0]), .i_data_2(C[92][0]), .o_data(mult_result_i[92][0]), .i_clk(i_clk));
Sub0000000002  u_00000002E3_Sub0000000002(.i_data_1(A[92][1]), .i_data_2(B[92][1]), .o_data(mult_result_r[92][1]), .i_clk(i_clk));
Sub0000000002  u_00000002E4_Sub0000000002(.i_data_1(B[92][1]), .i_data_2(C[92][1]), .o_data(mult_result_i[92][1]), .i_clk(i_clk));
Sub0000000002  u_00000002E5_Sub0000000002(.i_data_1(A[92][2]), .i_data_2(B[92][2]), .o_data(mult_result_r[92][2]), .i_clk(i_clk));
Sub0000000002  u_00000002E6_Sub0000000002(.i_data_1(B[92][2]), .i_data_2(C[92][2]), .o_data(mult_result_i[92][2]), .i_clk(i_clk));
Sub0000000002  u_00000002E7_Sub0000000002(.i_data_1(A[92][3]), .i_data_2(B[92][3]), .o_data(mult_result_r[92][3]), .i_clk(i_clk));
Sub0000000002  u_00000002E8_Sub0000000002(.i_data_1(B[92][3]), .i_data_2(C[92][3]), .o_data(mult_result_i[92][3]), .i_clk(i_clk));
Sub0000000002  u_00000002E9_Sub0000000002(.i_data_1(A[93][0]), .i_data_2(B[93][0]), .o_data(mult_result_r[93][0]), .i_clk(i_clk));
Sub0000000002  u_00000002EA_Sub0000000002(.i_data_1(B[93][0]), .i_data_2(C[93][0]), .o_data(mult_result_i[93][0]), .i_clk(i_clk));
Sub0000000002  u_00000002EB_Sub0000000002(.i_data_1(A[93][1]), .i_data_2(B[93][1]), .o_data(mult_result_r[93][1]), .i_clk(i_clk));
Sub0000000002  u_00000002EC_Sub0000000002(.i_data_1(B[93][1]), .i_data_2(C[93][1]), .o_data(mult_result_i[93][1]), .i_clk(i_clk));
Sub0000000002  u_00000002ED_Sub0000000002(.i_data_1(A[93][2]), .i_data_2(B[93][2]), .o_data(mult_result_r[93][2]), .i_clk(i_clk));
Sub0000000002  u_00000002EE_Sub0000000002(.i_data_1(B[93][2]), .i_data_2(C[93][2]), .o_data(mult_result_i[93][2]), .i_clk(i_clk));
Sub0000000002  u_00000002EF_Sub0000000002(.i_data_1(A[93][3]), .i_data_2(B[93][3]), .o_data(mult_result_r[93][3]), .i_clk(i_clk));
Sub0000000002  u_00000002F0_Sub0000000002(.i_data_1(B[93][3]), .i_data_2(C[93][3]), .o_data(mult_result_i[93][3]), .i_clk(i_clk));
Sub0000000002  u_00000002F1_Sub0000000002(.i_data_1(A[94][0]), .i_data_2(B[94][0]), .o_data(mult_result_r[94][0]), .i_clk(i_clk));
Sub0000000002  u_00000002F2_Sub0000000002(.i_data_1(B[94][0]), .i_data_2(C[94][0]), .o_data(mult_result_i[94][0]), .i_clk(i_clk));
Sub0000000002  u_00000002F3_Sub0000000002(.i_data_1(A[94][1]), .i_data_2(B[94][1]), .o_data(mult_result_r[94][1]), .i_clk(i_clk));
Sub0000000002  u_00000002F4_Sub0000000002(.i_data_1(B[94][1]), .i_data_2(C[94][1]), .o_data(mult_result_i[94][1]), .i_clk(i_clk));
Sub0000000002  u_00000002F5_Sub0000000002(.i_data_1(A[94][2]), .i_data_2(B[94][2]), .o_data(mult_result_r[94][2]), .i_clk(i_clk));
Sub0000000002  u_00000002F6_Sub0000000002(.i_data_1(B[94][2]), .i_data_2(C[94][2]), .o_data(mult_result_i[94][2]), .i_clk(i_clk));
Sub0000000002  u_00000002F7_Sub0000000002(.i_data_1(A[94][3]), .i_data_2(B[94][3]), .o_data(mult_result_r[94][3]), .i_clk(i_clk));
Sub0000000002  u_00000002F8_Sub0000000002(.i_data_1(B[94][3]), .i_data_2(C[94][3]), .o_data(mult_result_i[94][3]), .i_clk(i_clk));
Sub0000000002  u_00000002F9_Sub0000000002(.i_data_1(A[95][0]), .i_data_2(B[95][0]), .o_data(mult_result_r[95][0]), .i_clk(i_clk));
Sub0000000002  u_00000002FA_Sub0000000002(.i_data_1(B[95][0]), .i_data_2(C[95][0]), .o_data(mult_result_i[95][0]), .i_clk(i_clk));
Sub0000000002  u_00000002FB_Sub0000000002(.i_data_1(A[95][1]), .i_data_2(B[95][1]), .o_data(mult_result_r[95][1]), .i_clk(i_clk));
Sub0000000002  u_00000002FC_Sub0000000002(.i_data_1(B[95][1]), .i_data_2(C[95][1]), .o_data(mult_result_i[95][1]), .i_clk(i_clk));
Sub0000000002  u_00000002FD_Sub0000000002(.i_data_1(A[95][2]), .i_data_2(B[95][2]), .o_data(mult_result_r[95][2]), .i_clk(i_clk));
Sub0000000002  u_00000002FE_Sub0000000002(.i_data_1(B[95][2]), .i_data_2(C[95][2]), .o_data(mult_result_i[95][2]), .i_clk(i_clk));
Sub0000000002  u_00000002FF_Sub0000000002(.i_data_1(A[95][3]), .i_data_2(B[95][3]), .o_data(mult_result_r[95][3]), .i_clk(i_clk));
Sub0000000002  u_0000000300_Sub0000000002(.i_data_1(B[95][3]), .i_data_2(C[95][3]), .o_data(mult_result_i[95][3]), .i_clk(i_clk));
Sub0000000002  u_0000000301_Sub0000000002(.i_data_1(A[96][0]), .i_data_2(B[96][0]), .o_data(mult_result_r[96][0]), .i_clk(i_clk));
Sub0000000002  u_0000000302_Sub0000000002(.i_data_1(B[96][0]), .i_data_2(C[96][0]), .o_data(mult_result_i[96][0]), .i_clk(i_clk));
Sub0000000002  u_0000000303_Sub0000000002(.i_data_1(A[96][1]), .i_data_2(B[96][1]), .o_data(mult_result_r[96][1]), .i_clk(i_clk));
Sub0000000002  u_0000000304_Sub0000000002(.i_data_1(B[96][1]), .i_data_2(C[96][1]), .o_data(mult_result_i[96][1]), .i_clk(i_clk));
Sub0000000002  u_0000000305_Sub0000000002(.i_data_1(A[96][2]), .i_data_2(B[96][2]), .o_data(mult_result_r[96][2]), .i_clk(i_clk));
Sub0000000002  u_0000000306_Sub0000000002(.i_data_1(B[96][2]), .i_data_2(C[96][2]), .o_data(mult_result_i[96][2]), .i_clk(i_clk));
Sub0000000002  u_0000000307_Sub0000000002(.i_data_1(A[96][3]), .i_data_2(B[96][3]), .o_data(mult_result_r[96][3]), .i_clk(i_clk));
Sub0000000002  u_0000000308_Sub0000000002(.i_data_1(B[96][3]), .i_data_2(C[96][3]), .o_data(mult_result_i[96][3]), .i_clk(i_clk));
Sub0000000002  u_0000000309_Sub0000000002(.i_data_1(A[97][0]), .i_data_2(B[97][0]), .o_data(mult_result_r[97][0]), .i_clk(i_clk));
Sub0000000002  u_000000030A_Sub0000000002(.i_data_1(B[97][0]), .i_data_2(C[97][0]), .o_data(mult_result_i[97][0]), .i_clk(i_clk));
Sub0000000002  u_000000030B_Sub0000000002(.i_data_1(A[97][1]), .i_data_2(B[97][1]), .o_data(mult_result_r[97][1]), .i_clk(i_clk));
Sub0000000002  u_000000030C_Sub0000000002(.i_data_1(B[97][1]), .i_data_2(C[97][1]), .o_data(mult_result_i[97][1]), .i_clk(i_clk));
Sub0000000002  u_000000030D_Sub0000000002(.i_data_1(A[97][2]), .i_data_2(B[97][2]), .o_data(mult_result_r[97][2]), .i_clk(i_clk));
Sub0000000002  u_000000030E_Sub0000000002(.i_data_1(B[97][2]), .i_data_2(C[97][2]), .o_data(mult_result_i[97][2]), .i_clk(i_clk));
Sub0000000002  u_000000030F_Sub0000000002(.i_data_1(A[97][3]), .i_data_2(B[97][3]), .o_data(mult_result_r[97][3]), .i_clk(i_clk));
Sub0000000002  u_0000000310_Sub0000000002(.i_data_1(B[97][3]), .i_data_2(C[97][3]), .o_data(mult_result_i[97][3]), .i_clk(i_clk));
Sub0000000002  u_0000000311_Sub0000000002(.i_data_1(A[98][0]), .i_data_2(B[98][0]), .o_data(mult_result_r[98][0]), .i_clk(i_clk));
Sub0000000002  u_0000000312_Sub0000000002(.i_data_1(B[98][0]), .i_data_2(C[98][0]), .o_data(mult_result_i[98][0]), .i_clk(i_clk));
Sub0000000002  u_0000000313_Sub0000000002(.i_data_1(A[98][1]), .i_data_2(B[98][1]), .o_data(mult_result_r[98][1]), .i_clk(i_clk));
Sub0000000002  u_0000000314_Sub0000000002(.i_data_1(B[98][1]), .i_data_2(C[98][1]), .o_data(mult_result_i[98][1]), .i_clk(i_clk));
Sub0000000002  u_0000000315_Sub0000000002(.i_data_1(A[98][2]), .i_data_2(B[98][2]), .o_data(mult_result_r[98][2]), .i_clk(i_clk));
Sub0000000002  u_0000000316_Sub0000000002(.i_data_1(B[98][2]), .i_data_2(C[98][2]), .o_data(mult_result_i[98][2]), .i_clk(i_clk));
Sub0000000002  u_0000000317_Sub0000000002(.i_data_1(A[98][3]), .i_data_2(B[98][3]), .o_data(mult_result_r[98][3]), .i_clk(i_clk));
Sub0000000002  u_0000000318_Sub0000000002(.i_data_1(B[98][3]), .i_data_2(C[98][3]), .o_data(mult_result_i[98][3]), .i_clk(i_clk));
Sub0000000002  u_0000000319_Sub0000000002(.i_data_1(A[99][0]), .i_data_2(B[99][0]), .o_data(mult_result_r[99][0]), .i_clk(i_clk));
Sub0000000002  u_000000031A_Sub0000000002(.i_data_1(B[99][0]), .i_data_2(C[99][0]), .o_data(mult_result_i[99][0]), .i_clk(i_clk));
Sub0000000002  u_000000031B_Sub0000000002(.i_data_1(A[99][1]), .i_data_2(B[99][1]), .o_data(mult_result_r[99][1]), .i_clk(i_clk));
Sub0000000002  u_000000031C_Sub0000000002(.i_data_1(B[99][1]), .i_data_2(C[99][1]), .o_data(mult_result_i[99][1]), .i_clk(i_clk));
Sub0000000002  u_000000031D_Sub0000000002(.i_data_1(A[99][2]), .i_data_2(B[99][2]), .o_data(mult_result_r[99][2]), .i_clk(i_clk));
Sub0000000002  u_000000031E_Sub0000000002(.i_data_1(B[99][2]), .i_data_2(C[99][2]), .o_data(mult_result_i[99][2]), .i_clk(i_clk));
Sub0000000002  u_000000031F_Sub0000000002(.i_data_1(A[99][3]), .i_data_2(B[99][3]), .o_data(mult_result_r[99][3]), .i_clk(i_clk));
Sub0000000002  u_0000000320_Sub0000000002(.i_data_1(B[99][3]), .i_data_2(C[99][3]), .o_data(mult_result_i[99][3]), .i_clk(i_clk));
Sub0000000002  u_0000000321_Sub0000000002(.i_data_1(A[100][0]), .i_data_2(B[100][0]), .o_data(mult_result_r[100][0]), .i_clk(i_clk));
Sub0000000002  u_0000000322_Sub0000000002(.i_data_1(B[100][0]), .i_data_2(C[100][0]), .o_data(mult_result_i[100][0]), .i_clk(i_clk));
Sub0000000002  u_0000000323_Sub0000000002(.i_data_1(A[100][1]), .i_data_2(B[100][1]), .o_data(mult_result_r[100][1]), .i_clk(i_clk));
Sub0000000002  u_0000000324_Sub0000000002(.i_data_1(B[100][1]), .i_data_2(C[100][1]), .o_data(mult_result_i[100][1]), .i_clk(i_clk));
Sub0000000002  u_0000000325_Sub0000000002(.i_data_1(A[100][2]), .i_data_2(B[100][2]), .o_data(mult_result_r[100][2]), .i_clk(i_clk));
Sub0000000002  u_0000000326_Sub0000000002(.i_data_1(B[100][2]), .i_data_2(C[100][2]), .o_data(mult_result_i[100][2]), .i_clk(i_clk));
Sub0000000002  u_0000000327_Sub0000000002(.i_data_1(A[100][3]), .i_data_2(B[100][3]), .o_data(mult_result_r[100][3]), .i_clk(i_clk));
Sub0000000002  u_0000000328_Sub0000000002(.i_data_1(B[100][3]), .i_data_2(C[100][3]), .o_data(mult_result_i[100][3]), .i_clk(i_clk));
Sub0000000002  u_0000000329_Sub0000000002(.i_data_1(A[101][0]), .i_data_2(B[101][0]), .o_data(mult_result_r[101][0]), .i_clk(i_clk));
Sub0000000002  u_000000032A_Sub0000000002(.i_data_1(B[101][0]), .i_data_2(C[101][0]), .o_data(mult_result_i[101][0]), .i_clk(i_clk));
Sub0000000002  u_000000032B_Sub0000000002(.i_data_1(A[101][1]), .i_data_2(B[101][1]), .o_data(mult_result_r[101][1]), .i_clk(i_clk));
Sub0000000002  u_000000032C_Sub0000000002(.i_data_1(B[101][1]), .i_data_2(C[101][1]), .o_data(mult_result_i[101][1]), .i_clk(i_clk));
Sub0000000002  u_000000032D_Sub0000000002(.i_data_1(A[101][2]), .i_data_2(B[101][2]), .o_data(mult_result_r[101][2]), .i_clk(i_clk));
Sub0000000002  u_000000032E_Sub0000000002(.i_data_1(B[101][2]), .i_data_2(C[101][2]), .o_data(mult_result_i[101][2]), .i_clk(i_clk));
Sub0000000002  u_000000032F_Sub0000000002(.i_data_1(A[101][3]), .i_data_2(B[101][3]), .o_data(mult_result_r[101][3]), .i_clk(i_clk));
Sub0000000002  u_0000000330_Sub0000000002(.i_data_1(B[101][3]), .i_data_2(C[101][3]), .o_data(mult_result_i[101][3]), .i_clk(i_clk));
Sub0000000002  u_0000000331_Sub0000000002(.i_data_1(A[102][0]), .i_data_2(B[102][0]), .o_data(mult_result_r[102][0]), .i_clk(i_clk));
Sub0000000002  u_0000000332_Sub0000000002(.i_data_1(B[102][0]), .i_data_2(C[102][0]), .o_data(mult_result_i[102][0]), .i_clk(i_clk));
Sub0000000002  u_0000000333_Sub0000000002(.i_data_1(A[102][1]), .i_data_2(B[102][1]), .o_data(mult_result_r[102][1]), .i_clk(i_clk));
Sub0000000002  u_0000000334_Sub0000000002(.i_data_1(B[102][1]), .i_data_2(C[102][1]), .o_data(mult_result_i[102][1]), .i_clk(i_clk));
Sub0000000002  u_0000000335_Sub0000000002(.i_data_1(A[102][2]), .i_data_2(B[102][2]), .o_data(mult_result_r[102][2]), .i_clk(i_clk));
Sub0000000002  u_0000000336_Sub0000000002(.i_data_1(B[102][2]), .i_data_2(C[102][2]), .o_data(mult_result_i[102][2]), .i_clk(i_clk));
Sub0000000002  u_0000000337_Sub0000000002(.i_data_1(A[102][3]), .i_data_2(B[102][3]), .o_data(mult_result_r[102][3]), .i_clk(i_clk));
Sub0000000002  u_0000000338_Sub0000000002(.i_data_1(B[102][3]), .i_data_2(C[102][3]), .o_data(mult_result_i[102][3]), .i_clk(i_clk));
Sub0000000002  u_0000000339_Sub0000000002(.i_data_1(A[103][0]), .i_data_2(B[103][0]), .o_data(mult_result_r[103][0]), .i_clk(i_clk));
Sub0000000002  u_000000033A_Sub0000000002(.i_data_1(B[103][0]), .i_data_2(C[103][0]), .o_data(mult_result_i[103][0]), .i_clk(i_clk));
Sub0000000002  u_000000033B_Sub0000000002(.i_data_1(A[103][1]), .i_data_2(B[103][1]), .o_data(mult_result_r[103][1]), .i_clk(i_clk));
Sub0000000002  u_000000033C_Sub0000000002(.i_data_1(B[103][1]), .i_data_2(C[103][1]), .o_data(mult_result_i[103][1]), .i_clk(i_clk));
Sub0000000002  u_000000033D_Sub0000000002(.i_data_1(A[103][2]), .i_data_2(B[103][2]), .o_data(mult_result_r[103][2]), .i_clk(i_clk));
Sub0000000002  u_000000033E_Sub0000000002(.i_data_1(B[103][2]), .i_data_2(C[103][2]), .o_data(mult_result_i[103][2]), .i_clk(i_clk));
Sub0000000002  u_000000033F_Sub0000000002(.i_data_1(A[103][3]), .i_data_2(B[103][3]), .o_data(mult_result_r[103][3]), .i_clk(i_clk));
Sub0000000002  u_0000000340_Sub0000000002(.i_data_1(B[103][3]), .i_data_2(C[103][3]), .o_data(mult_result_i[103][3]), .i_clk(i_clk));
Sub0000000002  u_0000000341_Sub0000000002(.i_data_1(A[104][0]), .i_data_2(B[104][0]), .o_data(mult_result_r[104][0]), .i_clk(i_clk));
Sub0000000002  u_0000000342_Sub0000000002(.i_data_1(B[104][0]), .i_data_2(C[104][0]), .o_data(mult_result_i[104][0]), .i_clk(i_clk));
Sub0000000002  u_0000000343_Sub0000000002(.i_data_1(A[104][1]), .i_data_2(B[104][1]), .o_data(mult_result_r[104][1]), .i_clk(i_clk));
Sub0000000002  u_0000000344_Sub0000000002(.i_data_1(B[104][1]), .i_data_2(C[104][1]), .o_data(mult_result_i[104][1]), .i_clk(i_clk));
Sub0000000002  u_0000000345_Sub0000000002(.i_data_1(A[104][2]), .i_data_2(B[104][2]), .o_data(mult_result_r[104][2]), .i_clk(i_clk));
Sub0000000002  u_0000000346_Sub0000000002(.i_data_1(B[104][2]), .i_data_2(C[104][2]), .o_data(mult_result_i[104][2]), .i_clk(i_clk));
Sub0000000002  u_0000000347_Sub0000000002(.i_data_1(A[104][3]), .i_data_2(B[104][3]), .o_data(mult_result_r[104][3]), .i_clk(i_clk));
Sub0000000002  u_0000000348_Sub0000000002(.i_data_1(B[104][3]), .i_data_2(C[104][3]), .o_data(mult_result_i[104][3]), .i_clk(i_clk));
Sub0000000002  u_0000000349_Sub0000000002(.i_data_1(A[105][0]), .i_data_2(B[105][0]), .o_data(mult_result_r[105][0]), .i_clk(i_clk));
Sub0000000002  u_000000034A_Sub0000000002(.i_data_1(B[105][0]), .i_data_2(C[105][0]), .o_data(mult_result_i[105][0]), .i_clk(i_clk));
Sub0000000002  u_000000034B_Sub0000000002(.i_data_1(A[105][1]), .i_data_2(B[105][1]), .o_data(mult_result_r[105][1]), .i_clk(i_clk));
Sub0000000002  u_000000034C_Sub0000000002(.i_data_1(B[105][1]), .i_data_2(C[105][1]), .o_data(mult_result_i[105][1]), .i_clk(i_clk));
Sub0000000002  u_000000034D_Sub0000000002(.i_data_1(A[105][2]), .i_data_2(B[105][2]), .o_data(mult_result_r[105][2]), .i_clk(i_clk));
Sub0000000002  u_000000034E_Sub0000000002(.i_data_1(B[105][2]), .i_data_2(C[105][2]), .o_data(mult_result_i[105][2]), .i_clk(i_clk));
Sub0000000002  u_000000034F_Sub0000000002(.i_data_1(A[105][3]), .i_data_2(B[105][3]), .o_data(mult_result_r[105][3]), .i_clk(i_clk));
Sub0000000002  u_0000000350_Sub0000000002(.i_data_1(B[105][3]), .i_data_2(C[105][3]), .o_data(mult_result_i[105][3]), .i_clk(i_clk));
Sub0000000002  u_0000000351_Sub0000000002(.i_data_1(A[106][0]), .i_data_2(B[106][0]), .o_data(mult_result_r[106][0]), .i_clk(i_clk));
Sub0000000002  u_0000000352_Sub0000000002(.i_data_1(B[106][0]), .i_data_2(C[106][0]), .o_data(mult_result_i[106][0]), .i_clk(i_clk));
Sub0000000002  u_0000000353_Sub0000000002(.i_data_1(A[106][1]), .i_data_2(B[106][1]), .o_data(mult_result_r[106][1]), .i_clk(i_clk));
Sub0000000002  u_0000000354_Sub0000000002(.i_data_1(B[106][1]), .i_data_2(C[106][1]), .o_data(mult_result_i[106][1]), .i_clk(i_clk));
Sub0000000002  u_0000000355_Sub0000000002(.i_data_1(A[106][2]), .i_data_2(B[106][2]), .o_data(mult_result_r[106][2]), .i_clk(i_clk));
Sub0000000002  u_0000000356_Sub0000000002(.i_data_1(B[106][2]), .i_data_2(C[106][2]), .o_data(mult_result_i[106][2]), .i_clk(i_clk));
Sub0000000002  u_0000000357_Sub0000000002(.i_data_1(A[106][3]), .i_data_2(B[106][3]), .o_data(mult_result_r[106][3]), .i_clk(i_clk));
Sub0000000002  u_0000000358_Sub0000000002(.i_data_1(B[106][3]), .i_data_2(C[106][3]), .o_data(mult_result_i[106][3]), .i_clk(i_clk));
Sub0000000002  u_0000000359_Sub0000000002(.i_data_1(A[107][0]), .i_data_2(B[107][0]), .o_data(mult_result_r[107][0]), .i_clk(i_clk));
Sub0000000002  u_000000035A_Sub0000000002(.i_data_1(B[107][0]), .i_data_2(C[107][0]), .o_data(mult_result_i[107][0]), .i_clk(i_clk));
Sub0000000002  u_000000035B_Sub0000000002(.i_data_1(A[107][1]), .i_data_2(B[107][1]), .o_data(mult_result_r[107][1]), .i_clk(i_clk));
Sub0000000002  u_000000035C_Sub0000000002(.i_data_1(B[107][1]), .i_data_2(C[107][1]), .o_data(mult_result_i[107][1]), .i_clk(i_clk));
Sub0000000002  u_000000035D_Sub0000000002(.i_data_1(A[107][2]), .i_data_2(B[107][2]), .o_data(mult_result_r[107][2]), .i_clk(i_clk));
Sub0000000002  u_000000035E_Sub0000000002(.i_data_1(B[107][2]), .i_data_2(C[107][2]), .o_data(mult_result_i[107][2]), .i_clk(i_clk));
Sub0000000002  u_000000035F_Sub0000000002(.i_data_1(A[107][3]), .i_data_2(B[107][3]), .o_data(mult_result_r[107][3]), .i_clk(i_clk));
Sub0000000002  u_0000000360_Sub0000000002(.i_data_1(B[107][3]), .i_data_2(C[107][3]), .o_data(mult_result_i[107][3]), .i_clk(i_clk));
Sub0000000002  u_0000000361_Sub0000000002(.i_data_1(A[108][0]), .i_data_2(B[108][0]), .o_data(mult_result_r[108][0]), .i_clk(i_clk));
Sub0000000002  u_0000000362_Sub0000000002(.i_data_1(B[108][0]), .i_data_2(C[108][0]), .o_data(mult_result_i[108][0]), .i_clk(i_clk));
Sub0000000002  u_0000000363_Sub0000000002(.i_data_1(A[108][1]), .i_data_2(B[108][1]), .o_data(mult_result_r[108][1]), .i_clk(i_clk));
Sub0000000002  u_0000000364_Sub0000000002(.i_data_1(B[108][1]), .i_data_2(C[108][1]), .o_data(mult_result_i[108][1]), .i_clk(i_clk));
Sub0000000002  u_0000000365_Sub0000000002(.i_data_1(A[108][2]), .i_data_2(B[108][2]), .o_data(mult_result_r[108][2]), .i_clk(i_clk));
Sub0000000002  u_0000000366_Sub0000000002(.i_data_1(B[108][2]), .i_data_2(C[108][2]), .o_data(mult_result_i[108][2]), .i_clk(i_clk));
Sub0000000002  u_0000000367_Sub0000000002(.i_data_1(A[108][3]), .i_data_2(B[108][3]), .o_data(mult_result_r[108][3]), .i_clk(i_clk));
Sub0000000002  u_0000000368_Sub0000000002(.i_data_1(B[108][3]), .i_data_2(C[108][3]), .o_data(mult_result_i[108][3]), .i_clk(i_clk));
Sub0000000002  u_0000000369_Sub0000000002(.i_data_1(A[109][0]), .i_data_2(B[109][0]), .o_data(mult_result_r[109][0]), .i_clk(i_clk));
Sub0000000002  u_000000036A_Sub0000000002(.i_data_1(B[109][0]), .i_data_2(C[109][0]), .o_data(mult_result_i[109][0]), .i_clk(i_clk));
Sub0000000002  u_000000036B_Sub0000000002(.i_data_1(A[109][1]), .i_data_2(B[109][1]), .o_data(mult_result_r[109][1]), .i_clk(i_clk));
Sub0000000002  u_000000036C_Sub0000000002(.i_data_1(B[109][1]), .i_data_2(C[109][1]), .o_data(mult_result_i[109][1]), .i_clk(i_clk));
Sub0000000002  u_000000036D_Sub0000000002(.i_data_1(A[109][2]), .i_data_2(B[109][2]), .o_data(mult_result_r[109][2]), .i_clk(i_clk));
Sub0000000002  u_000000036E_Sub0000000002(.i_data_1(B[109][2]), .i_data_2(C[109][2]), .o_data(mult_result_i[109][2]), .i_clk(i_clk));
Sub0000000002  u_000000036F_Sub0000000002(.i_data_1(A[109][3]), .i_data_2(B[109][3]), .o_data(mult_result_r[109][3]), .i_clk(i_clk));
Sub0000000002  u_0000000370_Sub0000000002(.i_data_1(B[109][3]), .i_data_2(C[109][3]), .o_data(mult_result_i[109][3]), .i_clk(i_clk));
Sub0000000002  u_0000000371_Sub0000000002(.i_data_1(A[110][0]), .i_data_2(B[110][0]), .o_data(mult_result_r[110][0]), .i_clk(i_clk));
Sub0000000002  u_0000000372_Sub0000000002(.i_data_1(B[110][0]), .i_data_2(C[110][0]), .o_data(mult_result_i[110][0]), .i_clk(i_clk));
Sub0000000002  u_0000000373_Sub0000000002(.i_data_1(A[110][1]), .i_data_2(B[110][1]), .o_data(mult_result_r[110][1]), .i_clk(i_clk));
Sub0000000002  u_0000000374_Sub0000000002(.i_data_1(B[110][1]), .i_data_2(C[110][1]), .o_data(mult_result_i[110][1]), .i_clk(i_clk));
Sub0000000002  u_0000000375_Sub0000000002(.i_data_1(A[110][2]), .i_data_2(B[110][2]), .o_data(mult_result_r[110][2]), .i_clk(i_clk));
Sub0000000002  u_0000000376_Sub0000000002(.i_data_1(B[110][2]), .i_data_2(C[110][2]), .o_data(mult_result_i[110][2]), .i_clk(i_clk));
Sub0000000002  u_0000000377_Sub0000000002(.i_data_1(A[110][3]), .i_data_2(B[110][3]), .o_data(mult_result_r[110][3]), .i_clk(i_clk));
Sub0000000002  u_0000000378_Sub0000000002(.i_data_1(B[110][3]), .i_data_2(C[110][3]), .o_data(mult_result_i[110][3]), .i_clk(i_clk));
Sub0000000002  u_0000000379_Sub0000000002(.i_data_1(A[111][0]), .i_data_2(B[111][0]), .o_data(mult_result_r[111][0]), .i_clk(i_clk));
Sub0000000002  u_000000037A_Sub0000000002(.i_data_1(B[111][0]), .i_data_2(C[111][0]), .o_data(mult_result_i[111][0]), .i_clk(i_clk));
Sub0000000002  u_000000037B_Sub0000000002(.i_data_1(A[111][1]), .i_data_2(B[111][1]), .o_data(mult_result_r[111][1]), .i_clk(i_clk));
Sub0000000002  u_000000037C_Sub0000000002(.i_data_1(B[111][1]), .i_data_2(C[111][1]), .o_data(mult_result_i[111][1]), .i_clk(i_clk));
Sub0000000002  u_000000037D_Sub0000000002(.i_data_1(A[111][2]), .i_data_2(B[111][2]), .o_data(mult_result_r[111][2]), .i_clk(i_clk));
Sub0000000002  u_000000037E_Sub0000000002(.i_data_1(B[111][2]), .i_data_2(C[111][2]), .o_data(mult_result_i[111][2]), .i_clk(i_clk));
Sub0000000002  u_000000037F_Sub0000000002(.i_data_1(A[111][3]), .i_data_2(B[111][3]), .o_data(mult_result_r[111][3]), .i_clk(i_clk));
Sub0000000002  u_0000000380_Sub0000000002(.i_data_1(B[111][3]), .i_data_2(C[111][3]), .o_data(mult_result_i[111][3]), .i_clk(i_clk));
Sub0000000002  u_0000000381_Sub0000000002(.i_data_1(A[112][0]), .i_data_2(B[112][0]), .o_data(mult_result_r[112][0]), .i_clk(i_clk));
Sub0000000002  u_0000000382_Sub0000000002(.i_data_1(B[112][0]), .i_data_2(C[112][0]), .o_data(mult_result_i[112][0]), .i_clk(i_clk));
Sub0000000002  u_0000000383_Sub0000000002(.i_data_1(A[112][1]), .i_data_2(B[112][1]), .o_data(mult_result_r[112][1]), .i_clk(i_clk));
Sub0000000002  u_0000000384_Sub0000000002(.i_data_1(B[112][1]), .i_data_2(C[112][1]), .o_data(mult_result_i[112][1]), .i_clk(i_clk));
Sub0000000002  u_0000000385_Sub0000000002(.i_data_1(A[112][2]), .i_data_2(B[112][2]), .o_data(mult_result_r[112][2]), .i_clk(i_clk));
Sub0000000002  u_0000000386_Sub0000000002(.i_data_1(B[112][2]), .i_data_2(C[112][2]), .o_data(mult_result_i[112][2]), .i_clk(i_clk));
Sub0000000002  u_0000000387_Sub0000000002(.i_data_1(A[112][3]), .i_data_2(B[112][3]), .o_data(mult_result_r[112][3]), .i_clk(i_clk));
Sub0000000002  u_0000000388_Sub0000000002(.i_data_1(B[112][3]), .i_data_2(C[112][3]), .o_data(mult_result_i[112][3]), .i_clk(i_clk));
Sub0000000002  u_0000000389_Sub0000000002(.i_data_1(A[113][0]), .i_data_2(B[113][0]), .o_data(mult_result_r[113][0]), .i_clk(i_clk));
Sub0000000002  u_000000038A_Sub0000000002(.i_data_1(B[113][0]), .i_data_2(C[113][0]), .o_data(mult_result_i[113][0]), .i_clk(i_clk));
Sub0000000002  u_000000038B_Sub0000000002(.i_data_1(A[113][1]), .i_data_2(B[113][1]), .o_data(mult_result_r[113][1]), .i_clk(i_clk));
Sub0000000002  u_000000038C_Sub0000000002(.i_data_1(B[113][1]), .i_data_2(C[113][1]), .o_data(mult_result_i[113][1]), .i_clk(i_clk));
Sub0000000002  u_000000038D_Sub0000000002(.i_data_1(A[113][2]), .i_data_2(B[113][2]), .o_data(mult_result_r[113][2]), .i_clk(i_clk));
Sub0000000002  u_000000038E_Sub0000000002(.i_data_1(B[113][2]), .i_data_2(C[113][2]), .o_data(mult_result_i[113][2]), .i_clk(i_clk));
Sub0000000002  u_000000038F_Sub0000000002(.i_data_1(A[113][3]), .i_data_2(B[113][3]), .o_data(mult_result_r[113][3]), .i_clk(i_clk));
Sub0000000002  u_0000000390_Sub0000000002(.i_data_1(B[113][3]), .i_data_2(C[113][3]), .o_data(mult_result_i[113][3]), .i_clk(i_clk));
Sub0000000002  u_0000000391_Sub0000000002(.i_data_1(A[114][0]), .i_data_2(B[114][0]), .o_data(mult_result_r[114][0]), .i_clk(i_clk));
Sub0000000002  u_0000000392_Sub0000000002(.i_data_1(B[114][0]), .i_data_2(C[114][0]), .o_data(mult_result_i[114][0]), .i_clk(i_clk));
Sub0000000002  u_0000000393_Sub0000000002(.i_data_1(A[114][1]), .i_data_2(B[114][1]), .o_data(mult_result_r[114][1]), .i_clk(i_clk));
Sub0000000002  u_0000000394_Sub0000000002(.i_data_1(B[114][1]), .i_data_2(C[114][1]), .o_data(mult_result_i[114][1]), .i_clk(i_clk));
Sub0000000002  u_0000000395_Sub0000000002(.i_data_1(A[114][2]), .i_data_2(B[114][2]), .o_data(mult_result_r[114][2]), .i_clk(i_clk));
Sub0000000002  u_0000000396_Sub0000000002(.i_data_1(B[114][2]), .i_data_2(C[114][2]), .o_data(mult_result_i[114][2]), .i_clk(i_clk));
Sub0000000002  u_0000000397_Sub0000000002(.i_data_1(A[114][3]), .i_data_2(B[114][3]), .o_data(mult_result_r[114][3]), .i_clk(i_clk));
Sub0000000002  u_0000000398_Sub0000000002(.i_data_1(B[114][3]), .i_data_2(C[114][3]), .o_data(mult_result_i[114][3]), .i_clk(i_clk));
Sub0000000002  u_0000000399_Sub0000000002(.i_data_1(A[115][0]), .i_data_2(B[115][0]), .o_data(mult_result_r[115][0]), .i_clk(i_clk));
Sub0000000002  u_000000039A_Sub0000000002(.i_data_1(B[115][0]), .i_data_2(C[115][0]), .o_data(mult_result_i[115][0]), .i_clk(i_clk));
Sub0000000002  u_000000039B_Sub0000000002(.i_data_1(A[115][1]), .i_data_2(B[115][1]), .o_data(mult_result_r[115][1]), .i_clk(i_clk));
Sub0000000002  u_000000039C_Sub0000000002(.i_data_1(B[115][1]), .i_data_2(C[115][1]), .o_data(mult_result_i[115][1]), .i_clk(i_clk));
Sub0000000002  u_000000039D_Sub0000000002(.i_data_1(A[115][2]), .i_data_2(B[115][2]), .o_data(mult_result_r[115][2]), .i_clk(i_clk));
Sub0000000002  u_000000039E_Sub0000000002(.i_data_1(B[115][2]), .i_data_2(C[115][2]), .o_data(mult_result_i[115][2]), .i_clk(i_clk));
Sub0000000002  u_000000039F_Sub0000000002(.i_data_1(A[115][3]), .i_data_2(B[115][3]), .o_data(mult_result_r[115][3]), .i_clk(i_clk));
Sub0000000002  u_00000003A0_Sub0000000002(.i_data_1(B[115][3]), .i_data_2(C[115][3]), .o_data(mult_result_i[115][3]), .i_clk(i_clk));
Sub0000000002  u_00000003A1_Sub0000000002(.i_data_1(A[116][0]), .i_data_2(B[116][0]), .o_data(mult_result_r[116][0]), .i_clk(i_clk));
Sub0000000002  u_00000003A2_Sub0000000002(.i_data_1(B[116][0]), .i_data_2(C[116][0]), .o_data(mult_result_i[116][0]), .i_clk(i_clk));
Sub0000000002  u_00000003A3_Sub0000000002(.i_data_1(A[116][1]), .i_data_2(B[116][1]), .o_data(mult_result_r[116][1]), .i_clk(i_clk));
Sub0000000002  u_00000003A4_Sub0000000002(.i_data_1(B[116][1]), .i_data_2(C[116][1]), .o_data(mult_result_i[116][1]), .i_clk(i_clk));
Sub0000000002  u_00000003A5_Sub0000000002(.i_data_1(A[116][2]), .i_data_2(B[116][2]), .o_data(mult_result_r[116][2]), .i_clk(i_clk));
Sub0000000002  u_00000003A6_Sub0000000002(.i_data_1(B[116][2]), .i_data_2(C[116][2]), .o_data(mult_result_i[116][2]), .i_clk(i_clk));
Sub0000000002  u_00000003A7_Sub0000000002(.i_data_1(A[116][3]), .i_data_2(B[116][3]), .o_data(mult_result_r[116][3]), .i_clk(i_clk));
Sub0000000002  u_00000003A8_Sub0000000002(.i_data_1(B[116][3]), .i_data_2(C[116][3]), .o_data(mult_result_i[116][3]), .i_clk(i_clk));
Sub0000000002  u_00000003A9_Sub0000000002(.i_data_1(A[117][0]), .i_data_2(B[117][0]), .o_data(mult_result_r[117][0]), .i_clk(i_clk));
Sub0000000002  u_00000003AA_Sub0000000002(.i_data_1(B[117][0]), .i_data_2(C[117][0]), .o_data(mult_result_i[117][0]), .i_clk(i_clk));
Sub0000000002  u_00000003AB_Sub0000000002(.i_data_1(A[117][1]), .i_data_2(B[117][1]), .o_data(mult_result_r[117][1]), .i_clk(i_clk));
Sub0000000002  u_00000003AC_Sub0000000002(.i_data_1(B[117][1]), .i_data_2(C[117][1]), .o_data(mult_result_i[117][1]), .i_clk(i_clk));
Sub0000000002  u_00000003AD_Sub0000000002(.i_data_1(A[117][2]), .i_data_2(B[117][2]), .o_data(mult_result_r[117][2]), .i_clk(i_clk));
Sub0000000002  u_00000003AE_Sub0000000002(.i_data_1(B[117][2]), .i_data_2(C[117][2]), .o_data(mult_result_i[117][2]), .i_clk(i_clk));
Sub0000000002  u_00000003AF_Sub0000000002(.i_data_1(A[117][3]), .i_data_2(B[117][3]), .o_data(mult_result_r[117][3]), .i_clk(i_clk));
Sub0000000002  u_00000003B0_Sub0000000002(.i_data_1(B[117][3]), .i_data_2(C[117][3]), .o_data(mult_result_i[117][3]), .i_clk(i_clk));
Sub0000000002  u_00000003B1_Sub0000000002(.i_data_1(A[118][0]), .i_data_2(B[118][0]), .o_data(mult_result_r[118][0]), .i_clk(i_clk));
Sub0000000002  u_00000003B2_Sub0000000002(.i_data_1(B[118][0]), .i_data_2(C[118][0]), .o_data(mult_result_i[118][0]), .i_clk(i_clk));
Sub0000000002  u_00000003B3_Sub0000000002(.i_data_1(A[118][1]), .i_data_2(B[118][1]), .o_data(mult_result_r[118][1]), .i_clk(i_clk));
Sub0000000002  u_00000003B4_Sub0000000002(.i_data_1(B[118][1]), .i_data_2(C[118][1]), .o_data(mult_result_i[118][1]), .i_clk(i_clk));
Sub0000000002  u_00000003B5_Sub0000000002(.i_data_1(A[118][2]), .i_data_2(B[118][2]), .o_data(mult_result_r[118][2]), .i_clk(i_clk));
Sub0000000002  u_00000003B6_Sub0000000002(.i_data_1(B[118][2]), .i_data_2(C[118][2]), .o_data(mult_result_i[118][2]), .i_clk(i_clk));
Sub0000000002  u_00000003B7_Sub0000000002(.i_data_1(A[118][3]), .i_data_2(B[118][3]), .o_data(mult_result_r[118][3]), .i_clk(i_clk));
Sub0000000002  u_00000003B8_Sub0000000002(.i_data_1(B[118][3]), .i_data_2(C[118][3]), .o_data(mult_result_i[118][3]), .i_clk(i_clk));
Sub0000000002  u_00000003B9_Sub0000000002(.i_data_1(A[119][0]), .i_data_2(B[119][0]), .o_data(mult_result_r[119][0]), .i_clk(i_clk));
Sub0000000002  u_00000003BA_Sub0000000002(.i_data_1(B[119][0]), .i_data_2(C[119][0]), .o_data(mult_result_i[119][0]), .i_clk(i_clk));
Sub0000000002  u_00000003BB_Sub0000000002(.i_data_1(A[119][1]), .i_data_2(B[119][1]), .o_data(mult_result_r[119][1]), .i_clk(i_clk));
Sub0000000002  u_00000003BC_Sub0000000002(.i_data_1(B[119][1]), .i_data_2(C[119][1]), .o_data(mult_result_i[119][1]), .i_clk(i_clk));
Sub0000000002  u_00000003BD_Sub0000000002(.i_data_1(A[119][2]), .i_data_2(B[119][2]), .o_data(mult_result_r[119][2]), .i_clk(i_clk));
Sub0000000002  u_00000003BE_Sub0000000002(.i_data_1(B[119][2]), .i_data_2(C[119][2]), .o_data(mult_result_i[119][2]), .i_clk(i_clk));
Sub0000000002  u_00000003BF_Sub0000000002(.i_data_1(A[119][3]), .i_data_2(B[119][3]), .o_data(mult_result_r[119][3]), .i_clk(i_clk));
Sub0000000002  u_00000003C0_Sub0000000002(.i_data_1(B[119][3]), .i_data_2(C[119][3]), .o_data(mult_result_i[119][3]), .i_clk(i_clk));
Sub0000000002  u_00000003C1_Sub0000000002(.i_data_1(A[120][0]), .i_data_2(B[120][0]), .o_data(mult_result_r[120][0]), .i_clk(i_clk));
Sub0000000002  u_00000003C2_Sub0000000002(.i_data_1(B[120][0]), .i_data_2(C[120][0]), .o_data(mult_result_i[120][0]), .i_clk(i_clk));
Sub0000000002  u_00000003C3_Sub0000000002(.i_data_1(A[120][1]), .i_data_2(B[120][1]), .o_data(mult_result_r[120][1]), .i_clk(i_clk));
Sub0000000002  u_00000003C4_Sub0000000002(.i_data_1(B[120][1]), .i_data_2(C[120][1]), .o_data(mult_result_i[120][1]), .i_clk(i_clk));
Sub0000000002  u_00000003C5_Sub0000000002(.i_data_1(A[120][2]), .i_data_2(B[120][2]), .o_data(mult_result_r[120][2]), .i_clk(i_clk));
Sub0000000002  u_00000003C6_Sub0000000002(.i_data_1(B[120][2]), .i_data_2(C[120][2]), .o_data(mult_result_i[120][2]), .i_clk(i_clk));
Sub0000000002  u_00000003C7_Sub0000000002(.i_data_1(A[120][3]), .i_data_2(B[120][3]), .o_data(mult_result_r[120][3]), .i_clk(i_clk));
Sub0000000002  u_00000003C8_Sub0000000002(.i_data_1(B[120][3]), .i_data_2(C[120][3]), .o_data(mult_result_i[120][3]), .i_clk(i_clk));
Sub0000000002  u_00000003C9_Sub0000000002(.i_data_1(A[121][0]), .i_data_2(B[121][0]), .o_data(mult_result_r[121][0]), .i_clk(i_clk));
Sub0000000002  u_00000003CA_Sub0000000002(.i_data_1(B[121][0]), .i_data_2(C[121][0]), .o_data(mult_result_i[121][0]), .i_clk(i_clk));
Sub0000000002  u_00000003CB_Sub0000000002(.i_data_1(A[121][1]), .i_data_2(B[121][1]), .o_data(mult_result_r[121][1]), .i_clk(i_clk));
Sub0000000002  u_00000003CC_Sub0000000002(.i_data_1(B[121][1]), .i_data_2(C[121][1]), .o_data(mult_result_i[121][1]), .i_clk(i_clk));
Sub0000000002  u_00000003CD_Sub0000000002(.i_data_1(A[121][2]), .i_data_2(B[121][2]), .o_data(mult_result_r[121][2]), .i_clk(i_clk));
Sub0000000002  u_00000003CE_Sub0000000002(.i_data_1(B[121][2]), .i_data_2(C[121][2]), .o_data(mult_result_i[121][2]), .i_clk(i_clk));
Sub0000000002  u_00000003CF_Sub0000000002(.i_data_1(A[121][3]), .i_data_2(B[121][3]), .o_data(mult_result_r[121][3]), .i_clk(i_clk));
Sub0000000002  u_00000003D0_Sub0000000002(.i_data_1(B[121][3]), .i_data_2(C[121][3]), .o_data(mult_result_i[121][3]), .i_clk(i_clk));
Sub0000000002  u_00000003D1_Sub0000000002(.i_data_1(A[122][0]), .i_data_2(B[122][0]), .o_data(mult_result_r[122][0]), .i_clk(i_clk));
Sub0000000002  u_00000003D2_Sub0000000002(.i_data_1(B[122][0]), .i_data_2(C[122][0]), .o_data(mult_result_i[122][0]), .i_clk(i_clk));
Sub0000000002  u_00000003D3_Sub0000000002(.i_data_1(A[122][1]), .i_data_2(B[122][1]), .o_data(mult_result_r[122][1]), .i_clk(i_clk));
Sub0000000002  u_00000003D4_Sub0000000002(.i_data_1(B[122][1]), .i_data_2(C[122][1]), .o_data(mult_result_i[122][1]), .i_clk(i_clk));
Sub0000000002  u_00000003D5_Sub0000000002(.i_data_1(A[122][2]), .i_data_2(B[122][2]), .o_data(mult_result_r[122][2]), .i_clk(i_clk));
Sub0000000002  u_00000003D6_Sub0000000002(.i_data_1(B[122][2]), .i_data_2(C[122][2]), .o_data(mult_result_i[122][2]), .i_clk(i_clk));
Sub0000000002  u_00000003D7_Sub0000000002(.i_data_1(A[122][3]), .i_data_2(B[122][3]), .o_data(mult_result_r[122][3]), .i_clk(i_clk));
Sub0000000002  u_00000003D8_Sub0000000002(.i_data_1(B[122][3]), .i_data_2(C[122][3]), .o_data(mult_result_i[122][3]), .i_clk(i_clk));
Sub0000000002  u_00000003D9_Sub0000000002(.i_data_1(A[123][0]), .i_data_2(B[123][0]), .o_data(mult_result_r[123][0]), .i_clk(i_clk));
Sub0000000002  u_00000003DA_Sub0000000002(.i_data_1(B[123][0]), .i_data_2(C[123][0]), .o_data(mult_result_i[123][0]), .i_clk(i_clk));
Sub0000000002  u_00000003DB_Sub0000000002(.i_data_1(A[123][1]), .i_data_2(B[123][1]), .o_data(mult_result_r[123][1]), .i_clk(i_clk));
Sub0000000002  u_00000003DC_Sub0000000002(.i_data_1(B[123][1]), .i_data_2(C[123][1]), .o_data(mult_result_i[123][1]), .i_clk(i_clk));
Sub0000000002  u_00000003DD_Sub0000000002(.i_data_1(A[123][2]), .i_data_2(B[123][2]), .o_data(mult_result_r[123][2]), .i_clk(i_clk));
Sub0000000002  u_00000003DE_Sub0000000002(.i_data_1(B[123][2]), .i_data_2(C[123][2]), .o_data(mult_result_i[123][2]), .i_clk(i_clk));
Sub0000000002  u_00000003DF_Sub0000000002(.i_data_1(A[123][3]), .i_data_2(B[123][3]), .o_data(mult_result_r[123][3]), .i_clk(i_clk));
Sub0000000002  u_00000003E0_Sub0000000002(.i_data_1(B[123][3]), .i_data_2(C[123][3]), .o_data(mult_result_i[123][3]), .i_clk(i_clk));
Sub0000000002  u_00000003E1_Sub0000000002(.i_data_1(A[124][0]), .i_data_2(B[124][0]), .o_data(mult_result_r[124][0]), .i_clk(i_clk));
Sub0000000002  u_00000003E2_Sub0000000002(.i_data_1(B[124][0]), .i_data_2(C[124][0]), .o_data(mult_result_i[124][0]), .i_clk(i_clk));
Sub0000000002  u_00000003E3_Sub0000000002(.i_data_1(A[124][1]), .i_data_2(B[124][1]), .o_data(mult_result_r[124][1]), .i_clk(i_clk));
Sub0000000002  u_00000003E4_Sub0000000002(.i_data_1(B[124][1]), .i_data_2(C[124][1]), .o_data(mult_result_i[124][1]), .i_clk(i_clk));
Sub0000000002  u_00000003E5_Sub0000000002(.i_data_1(A[124][2]), .i_data_2(B[124][2]), .o_data(mult_result_r[124][2]), .i_clk(i_clk));
Sub0000000002  u_00000003E6_Sub0000000002(.i_data_1(B[124][2]), .i_data_2(C[124][2]), .o_data(mult_result_i[124][2]), .i_clk(i_clk));
Sub0000000002  u_00000003E7_Sub0000000002(.i_data_1(A[124][3]), .i_data_2(B[124][3]), .o_data(mult_result_r[124][3]), .i_clk(i_clk));
Sub0000000002  u_00000003E8_Sub0000000002(.i_data_1(B[124][3]), .i_data_2(C[124][3]), .o_data(mult_result_i[124][3]), .i_clk(i_clk));
Sub0000000002  u_00000003E9_Sub0000000002(.i_data_1(A[125][0]), .i_data_2(B[125][0]), .o_data(mult_result_r[125][0]), .i_clk(i_clk));
Sub0000000002  u_00000003EA_Sub0000000002(.i_data_1(B[125][0]), .i_data_2(C[125][0]), .o_data(mult_result_i[125][0]), .i_clk(i_clk));
Sub0000000002  u_00000003EB_Sub0000000002(.i_data_1(A[125][1]), .i_data_2(B[125][1]), .o_data(mult_result_r[125][1]), .i_clk(i_clk));
Sub0000000002  u_00000003EC_Sub0000000002(.i_data_1(B[125][1]), .i_data_2(C[125][1]), .o_data(mult_result_i[125][1]), .i_clk(i_clk));
Sub0000000002  u_00000003ED_Sub0000000002(.i_data_1(A[125][2]), .i_data_2(B[125][2]), .o_data(mult_result_r[125][2]), .i_clk(i_clk));
Sub0000000002  u_00000003EE_Sub0000000002(.i_data_1(B[125][2]), .i_data_2(C[125][2]), .o_data(mult_result_i[125][2]), .i_clk(i_clk));
Sub0000000002  u_00000003EF_Sub0000000002(.i_data_1(A[125][3]), .i_data_2(B[125][3]), .o_data(mult_result_r[125][3]), .i_clk(i_clk));
Sub0000000002  u_00000003F0_Sub0000000002(.i_data_1(B[125][3]), .i_data_2(C[125][3]), .o_data(mult_result_i[125][3]), .i_clk(i_clk));
Sub0000000002  u_00000003F1_Sub0000000002(.i_data_1(A[126][0]), .i_data_2(B[126][0]), .o_data(mult_result_r[126][0]), .i_clk(i_clk));
Sub0000000002  u_00000003F2_Sub0000000002(.i_data_1(B[126][0]), .i_data_2(C[126][0]), .o_data(mult_result_i[126][0]), .i_clk(i_clk));
Sub0000000002  u_00000003F3_Sub0000000002(.i_data_1(A[126][1]), .i_data_2(B[126][1]), .o_data(mult_result_r[126][1]), .i_clk(i_clk));
Sub0000000002  u_00000003F4_Sub0000000002(.i_data_1(B[126][1]), .i_data_2(C[126][1]), .o_data(mult_result_i[126][1]), .i_clk(i_clk));
Sub0000000002  u_00000003F5_Sub0000000002(.i_data_1(A[126][2]), .i_data_2(B[126][2]), .o_data(mult_result_r[126][2]), .i_clk(i_clk));
Sub0000000002  u_00000003F6_Sub0000000002(.i_data_1(B[126][2]), .i_data_2(C[126][2]), .o_data(mult_result_i[126][2]), .i_clk(i_clk));
Sub0000000002  u_00000003F7_Sub0000000002(.i_data_1(A[126][3]), .i_data_2(B[126][3]), .o_data(mult_result_r[126][3]), .i_clk(i_clk));
Sub0000000002  u_00000003F8_Sub0000000002(.i_data_1(B[126][3]), .i_data_2(C[126][3]), .o_data(mult_result_i[126][3]), .i_clk(i_clk));
Sub0000000002  u_00000003F9_Sub0000000002(.i_data_1(A[127][0]), .i_data_2(B[127][0]), .o_data(mult_result_r[127][0]), .i_clk(i_clk));
Sub0000000002  u_00000003FA_Sub0000000002(.i_data_1(B[127][0]), .i_data_2(C[127][0]), .o_data(mult_result_i[127][0]), .i_clk(i_clk));
Sub0000000002  u_00000003FB_Sub0000000002(.i_data_1(A[127][1]), .i_data_2(B[127][1]), .o_data(mult_result_r[127][1]), .i_clk(i_clk));
Sub0000000002  u_00000003FC_Sub0000000002(.i_data_1(B[127][1]), .i_data_2(C[127][1]), .o_data(mult_result_i[127][1]), .i_clk(i_clk));
Sub0000000002  u_00000003FD_Sub0000000002(.i_data_1(A[127][2]), .i_data_2(B[127][2]), .o_data(mult_result_r[127][2]), .i_clk(i_clk));
Sub0000000002  u_00000003FE_Sub0000000002(.i_data_1(B[127][2]), .i_data_2(C[127][2]), .o_data(mult_result_i[127][2]), .i_clk(i_clk));
Sub0000000002  u_00000003FF_Sub0000000002(.i_data_1(A[127][3]), .i_data_2(B[127][3]), .o_data(mult_result_r[127][3]), .i_clk(i_clk));
Sub0000000002  u_0000000400_Sub0000000002(.i_data_1(B[127][3]), .i_data_2(C[127][3]), .o_data(mult_result_i[127][3]), .i_clk(i_clk));
Sub0000000002  u_0000000401_Sub0000000002(.i_data_1(A[128][0]), .i_data_2(B[128][0]), .o_data(mult_result_r[128][0]), .i_clk(i_clk));
Sub0000000002  u_0000000402_Sub0000000002(.i_data_1(B[128][0]), .i_data_2(C[128][0]), .o_data(mult_result_i[128][0]), .i_clk(i_clk));
Sub0000000002  u_0000000403_Sub0000000002(.i_data_1(A[128][1]), .i_data_2(B[128][1]), .o_data(mult_result_r[128][1]), .i_clk(i_clk));
Sub0000000002  u_0000000404_Sub0000000002(.i_data_1(B[128][1]), .i_data_2(C[128][1]), .o_data(mult_result_i[128][1]), .i_clk(i_clk));
Sub0000000002  u_0000000405_Sub0000000002(.i_data_1(A[128][2]), .i_data_2(B[128][2]), .o_data(mult_result_r[128][2]), .i_clk(i_clk));
Sub0000000002  u_0000000406_Sub0000000002(.i_data_1(B[128][2]), .i_data_2(C[128][2]), .o_data(mult_result_i[128][2]), .i_clk(i_clk));
Sub0000000002  u_0000000407_Sub0000000002(.i_data_1(A[128][3]), .i_data_2(B[128][3]), .o_data(mult_result_r[128][3]), .i_clk(i_clk));
Sub0000000002  u_0000000408_Sub0000000002(.i_data_1(B[128][3]), .i_data_2(C[128][3]), .o_data(mult_result_i[128][3]), .i_clk(i_clk));
Sub0000000002  u_0000000409_Sub0000000002(.i_data_1(A[129][0]), .i_data_2(B[129][0]), .o_data(mult_result_r[129][0]), .i_clk(i_clk));
Sub0000000002  u_000000040A_Sub0000000002(.i_data_1(B[129][0]), .i_data_2(C[129][0]), .o_data(mult_result_i[129][0]), .i_clk(i_clk));
Sub0000000002  u_000000040B_Sub0000000002(.i_data_1(A[129][1]), .i_data_2(B[129][1]), .o_data(mult_result_r[129][1]), .i_clk(i_clk));
Sub0000000002  u_000000040C_Sub0000000002(.i_data_1(B[129][1]), .i_data_2(C[129][1]), .o_data(mult_result_i[129][1]), .i_clk(i_clk));
Sub0000000002  u_000000040D_Sub0000000002(.i_data_1(A[129][2]), .i_data_2(B[129][2]), .o_data(mult_result_r[129][2]), .i_clk(i_clk));
Sub0000000002  u_000000040E_Sub0000000002(.i_data_1(B[129][2]), .i_data_2(C[129][2]), .o_data(mult_result_i[129][2]), .i_clk(i_clk));
Sub0000000002  u_000000040F_Sub0000000002(.i_data_1(A[129][3]), .i_data_2(B[129][3]), .o_data(mult_result_r[129][3]), .i_clk(i_clk));
Sub0000000002  u_0000000410_Sub0000000002(.i_data_1(B[129][3]), .i_data_2(C[129][3]), .o_data(mult_result_i[129][3]), .i_clk(i_clk));
Sub0000000002  u_0000000411_Sub0000000002(.i_data_1(A[130][0]), .i_data_2(B[130][0]), .o_data(mult_result_r[130][0]), .i_clk(i_clk));
Sub0000000002  u_0000000412_Sub0000000002(.i_data_1(B[130][0]), .i_data_2(C[130][0]), .o_data(mult_result_i[130][0]), .i_clk(i_clk));
Sub0000000002  u_0000000413_Sub0000000002(.i_data_1(A[130][1]), .i_data_2(B[130][1]), .o_data(mult_result_r[130][1]), .i_clk(i_clk));
Sub0000000002  u_0000000414_Sub0000000002(.i_data_1(B[130][1]), .i_data_2(C[130][1]), .o_data(mult_result_i[130][1]), .i_clk(i_clk));
Sub0000000002  u_0000000415_Sub0000000002(.i_data_1(A[130][2]), .i_data_2(B[130][2]), .o_data(mult_result_r[130][2]), .i_clk(i_clk));
Sub0000000002  u_0000000416_Sub0000000002(.i_data_1(B[130][2]), .i_data_2(C[130][2]), .o_data(mult_result_i[130][2]), .i_clk(i_clk));
Sub0000000002  u_0000000417_Sub0000000002(.i_data_1(A[130][3]), .i_data_2(B[130][3]), .o_data(mult_result_r[130][3]), .i_clk(i_clk));
Sub0000000002  u_0000000418_Sub0000000002(.i_data_1(B[130][3]), .i_data_2(C[130][3]), .o_data(mult_result_i[130][3]), .i_clk(i_clk));
Sub0000000002  u_0000000419_Sub0000000002(.i_data_1(A[131][0]), .i_data_2(B[131][0]), .o_data(mult_result_r[131][0]), .i_clk(i_clk));
Sub0000000002  u_000000041A_Sub0000000002(.i_data_1(B[131][0]), .i_data_2(C[131][0]), .o_data(mult_result_i[131][0]), .i_clk(i_clk));
Sub0000000002  u_000000041B_Sub0000000002(.i_data_1(A[131][1]), .i_data_2(B[131][1]), .o_data(mult_result_r[131][1]), .i_clk(i_clk));
Sub0000000002  u_000000041C_Sub0000000002(.i_data_1(B[131][1]), .i_data_2(C[131][1]), .o_data(mult_result_i[131][1]), .i_clk(i_clk));
Sub0000000002  u_000000041D_Sub0000000002(.i_data_1(A[131][2]), .i_data_2(B[131][2]), .o_data(mult_result_r[131][2]), .i_clk(i_clk));
Sub0000000002  u_000000041E_Sub0000000002(.i_data_1(B[131][2]), .i_data_2(C[131][2]), .o_data(mult_result_i[131][2]), .i_clk(i_clk));
Sub0000000002  u_000000041F_Sub0000000002(.i_data_1(A[131][3]), .i_data_2(B[131][3]), .o_data(mult_result_r[131][3]), .i_clk(i_clk));
Sub0000000002  u_0000000420_Sub0000000002(.i_data_1(B[131][3]), .i_data_2(C[131][3]), .o_data(mult_result_i[131][3]), .i_clk(i_clk));
Sub0000000002  u_0000000421_Sub0000000002(.i_data_1(A[132][0]), .i_data_2(B[132][0]), .o_data(mult_result_r[132][0]), .i_clk(i_clk));
Sub0000000002  u_0000000422_Sub0000000002(.i_data_1(B[132][0]), .i_data_2(C[132][0]), .o_data(mult_result_i[132][0]), .i_clk(i_clk));
Sub0000000002  u_0000000423_Sub0000000002(.i_data_1(A[132][1]), .i_data_2(B[132][1]), .o_data(mult_result_r[132][1]), .i_clk(i_clk));
Sub0000000002  u_0000000424_Sub0000000002(.i_data_1(B[132][1]), .i_data_2(C[132][1]), .o_data(mult_result_i[132][1]), .i_clk(i_clk));
Sub0000000002  u_0000000425_Sub0000000002(.i_data_1(A[132][2]), .i_data_2(B[132][2]), .o_data(mult_result_r[132][2]), .i_clk(i_clk));
Sub0000000002  u_0000000426_Sub0000000002(.i_data_1(B[132][2]), .i_data_2(C[132][2]), .o_data(mult_result_i[132][2]), .i_clk(i_clk));
Sub0000000002  u_0000000427_Sub0000000002(.i_data_1(A[132][3]), .i_data_2(B[132][3]), .o_data(mult_result_r[132][3]), .i_clk(i_clk));
Sub0000000002  u_0000000428_Sub0000000002(.i_data_1(B[132][3]), .i_data_2(C[132][3]), .o_data(mult_result_i[132][3]), .i_clk(i_clk));
Sub0000000002  u_0000000429_Sub0000000002(.i_data_1(A[133][0]), .i_data_2(B[133][0]), .o_data(mult_result_r[133][0]), .i_clk(i_clk));
Sub0000000002  u_000000042A_Sub0000000002(.i_data_1(B[133][0]), .i_data_2(C[133][0]), .o_data(mult_result_i[133][0]), .i_clk(i_clk));
Sub0000000002  u_000000042B_Sub0000000002(.i_data_1(A[133][1]), .i_data_2(B[133][1]), .o_data(mult_result_r[133][1]), .i_clk(i_clk));
Sub0000000002  u_000000042C_Sub0000000002(.i_data_1(B[133][1]), .i_data_2(C[133][1]), .o_data(mult_result_i[133][1]), .i_clk(i_clk));
Sub0000000002  u_000000042D_Sub0000000002(.i_data_1(A[133][2]), .i_data_2(B[133][2]), .o_data(mult_result_r[133][2]), .i_clk(i_clk));
Sub0000000002  u_000000042E_Sub0000000002(.i_data_1(B[133][2]), .i_data_2(C[133][2]), .o_data(mult_result_i[133][2]), .i_clk(i_clk));
Sub0000000002  u_000000042F_Sub0000000002(.i_data_1(A[133][3]), .i_data_2(B[133][3]), .o_data(mult_result_r[133][3]), .i_clk(i_clk));
Sub0000000002  u_0000000430_Sub0000000002(.i_data_1(B[133][3]), .i_data_2(C[133][3]), .o_data(mult_result_i[133][3]), .i_clk(i_clk));
Sub0000000002  u_0000000431_Sub0000000002(.i_data_1(A[134][0]), .i_data_2(B[134][0]), .o_data(mult_result_r[134][0]), .i_clk(i_clk));
Sub0000000002  u_0000000432_Sub0000000002(.i_data_1(B[134][0]), .i_data_2(C[134][0]), .o_data(mult_result_i[134][0]), .i_clk(i_clk));
Sub0000000002  u_0000000433_Sub0000000002(.i_data_1(A[134][1]), .i_data_2(B[134][1]), .o_data(mult_result_r[134][1]), .i_clk(i_clk));
Sub0000000002  u_0000000434_Sub0000000002(.i_data_1(B[134][1]), .i_data_2(C[134][1]), .o_data(mult_result_i[134][1]), .i_clk(i_clk));
Sub0000000002  u_0000000435_Sub0000000002(.i_data_1(A[134][2]), .i_data_2(B[134][2]), .o_data(mult_result_r[134][2]), .i_clk(i_clk));
Sub0000000002  u_0000000436_Sub0000000002(.i_data_1(B[134][2]), .i_data_2(C[134][2]), .o_data(mult_result_i[134][2]), .i_clk(i_clk));
Sub0000000002  u_0000000437_Sub0000000002(.i_data_1(A[134][3]), .i_data_2(B[134][3]), .o_data(mult_result_r[134][3]), .i_clk(i_clk));
Sub0000000002  u_0000000438_Sub0000000002(.i_data_1(B[134][3]), .i_data_2(C[134][3]), .o_data(mult_result_i[134][3]), .i_clk(i_clk));
Sub0000000002  u_0000000439_Sub0000000002(.i_data_1(A[135][0]), .i_data_2(B[135][0]), .o_data(mult_result_r[135][0]), .i_clk(i_clk));
Sub0000000002  u_000000043A_Sub0000000002(.i_data_1(B[135][0]), .i_data_2(C[135][0]), .o_data(mult_result_i[135][0]), .i_clk(i_clk));
Sub0000000002  u_000000043B_Sub0000000002(.i_data_1(A[135][1]), .i_data_2(B[135][1]), .o_data(mult_result_r[135][1]), .i_clk(i_clk));
Sub0000000002  u_000000043C_Sub0000000002(.i_data_1(B[135][1]), .i_data_2(C[135][1]), .o_data(mult_result_i[135][1]), .i_clk(i_clk));
Sub0000000002  u_000000043D_Sub0000000002(.i_data_1(A[135][2]), .i_data_2(B[135][2]), .o_data(mult_result_r[135][2]), .i_clk(i_clk));
Sub0000000002  u_000000043E_Sub0000000002(.i_data_1(B[135][2]), .i_data_2(C[135][2]), .o_data(mult_result_i[135][2]), .i_clk(i_clk));
Sub0000000002  u_000000043F_Sub0000000002(.i_data_1(A[135][3]), .i_data_2(B[135][3]), .o_data(mult_result_r[135][3]), .i_clk(i_clk));
Sub0000000002  u_0000000440_Sub0000000002(.i_data_1(B[135][3]), .i_data_2(C[135][3]), .o_data(mult_result_i[135][3]), .i_clk(i_clk));
Sub0000000002  u_0000000441_Sub0000000002(.i_data_1(A[136][0]), .i_data_2(B[136][0]), .o_data(mult_result_r[136][0]), .i_clk(i_clk));
Sub0000000002  u_0000000442_Sub0000000002(.i_data_1(B[136][0]), .i_data_2(C[136][0]), .o_data(mult_result_i[136][0]), .i_clk(i_clk));
Sub0000000002  u_0000000443_Sub0000000002(.i_data_1(A[136][1]), .i_data_2(B[136][1]), .o_data(mult_result_r[136][1]), .i_clk(i_clk));
Sub0000000002  u_0000000444_Sub0000000002(.i_data_1(B[136][1]), .i_data_2(C[136][1]), .o_data(mult_result_i[136][1]), .i_clk(i_clk));
Sub0000000002  u_0000000445_Sub0000000002(.i_data_1(A[136][2]), .i_data_2(B[136][2]), .o_data(mult_result_r[136][2]), .i_clk(i_clk));
Sub0000000002  u_0000000446_Sub0000000002(.i_data_1(B[136][2]), .i_data_2(C[136][2]), .o_data(mult_result_i[136][2]), .i_clk(i_clk));
Sub0000000002  u_0000000447_Sub0000000002(.i_data_1(A[136][3]), .i_data_2(B[136][3]), .o_data(mult_result_r[136][3]), .i_clk(i_clk));
Sub0000000002  u_0000000448_Sub0000000002(.i_data_1(B[136][3]), .i_data_2(C[136][3]), .o_data(mult_result_i[136][3]), .i_clk(i_clk));
Sub0000000002  u_0000000449_Sub0000000002(.i_data_1(A[137][0]), .i_data_2(B[137][0]), .o_data(mult_result_r[137][0]), .i_clk(i_clk));
Sub0000000002  u_000000044A_Sub0000000002(.i_data_1(B[137][0]), .i_data_2(C[137][0]), .o_data(mult_result_i[137][0]), .i_clk(i_clk));
Sub0000000002  u_000000044B_Sub0000000002(.i_data_1(A[137][1]), .i_data_2(B[137][1]), .o_data(mult_result_r[137][1]), .i_clk(i_clk));
Sub0000000002  u_000000044C_Sub0000000002(.i_data_1(B[137][1]), .i_data_2(C[137][1]), .o_data(mult_result_i[137][1]), .i_clk(i_clk));
Sub0000000002  u_000000044D_Sub0000000002(.i_data_1(A[137][2]), .i_data_2(B[137][2]), .o_data(mult_result_r[137][2]), .i_clk(i_clk));
Sub0000000002  u_000000044E_Sub0000000002(.i_data_1(B[137][2]), .i_data_2(C[137][2]), .o_data(mult_result_i[137][2]), .i_clk(i_clk));
Sub0000000002  u_000000044F_Sub0000000002(.i_data_1(A[137][3]), .i_data_2(B[137][3]), .o_data(mult_result_r[137][3]), .i_clk(i_clk));
Sub0000000002  u_0000000450_Sub0000000002(.i_data_1(B[137][3]), .i_data_2(C[137][3]), .o_data(mult_result_i[137][3]), .i_clk(i_clk));
Sub0000000002  u_0000000451_Sub0000000002(.i_data_1(A[138][0]), .i_data_2(B[138][0]), .o_data(mult_result_r[138][0]), .i_clk(i_clk));
Sub0000000002  u_0000000452_Sub0000000002(.i_data_1(B[138][0]), .i_data_2(C[138][0]), .o_data(mult_result_i[138][0]), .i_clk(i_clk));
Sub0000000002  u_0000000453_Sub0000000002(.i_data_1(A[138][1]), .i_data_2(B[138][1]), .o_data(mult_result_r[138][1]), .i_clk(i_clk));
Sub0000000002  u_0000000454_Sub0000000002(.i_data_1(B[138][1]), .i_data_2(C[138][1]), .o_data(mult_result_i[138][1]), .i_clk(i_clk));
Sub0000000002  u_0000000455_Sub0000000002(.i_data_1(A[138][2]), .i_data_2(B[138][2]), .o_data(mult_result_r[138][2]), .i_clk(i_clk));
Sub0000000002  u_0000000456_Sub0000000002(.i_data_1(B[138][2]), .i_data_2(C[138][2]), .o_data(mult_result_i[138][2]), .i_clk(i_clk));
Sub0000000002  u_0000000457_Sub0000000002(.i_data_1(A[138][3]), .i_data_2(B[138][3]), .o_data(mult_result_r[138][3]), .i_clk(i_clk));
Sub0000000002  u_0000000458_Sub0000000002(.i_data_1(B[138][3]), .i_data_2(C[138][3]), .o_data(mult_result_i[138][3]), .i_clk(i_clk));
Sub0000000002  u_0000000459_Sub0000000002(.i_data_1(A[139][0]), .i_data_2(B[139][0]), .o_data(mult_result_r[139][0]), .i_clk(i_clk));
Sub0000000002  u_000000045A_Sub0000000002(.i_data_1(B[139][0]), .i_data_2(C[139][0]), .o_data(mult_result_i[139][0]), .i_clk(i_clk));
Sub0000000002  u_000000045B_Sub0000000002(.i_data_1(A[139][1]), .i_data_2(B[139][1]), .o_data(mult_result_r[139][1]), .i_clk(i_clk));
Sub0000000002  u_000000045C_Sub0000000002(.i_data_1(B[139][1]), .i_data_2(C[139][1]), .o_data(mult_result_i[139][1]), .i_clk(i_clk));
Sub0000000002  u_000000045D_Sub0000000002(.i_data_1(A[139][2]), .i_data_2(B[139][2]), .o_data(mult_result_r[139][2]), .i_clk(i_clk));
Sub0000000002  u_000000045E_Sub0000000002(.i_data_1(B[139][2]), .i_data_2(C[139][2]), .o_data(mult_result_i[139][2]), .i_clk(i_clk));
Sub0000000002  u_000000045F_Sub0000000002(.i_data_1(A[139][3]), .i_data_2(B[139][3]), .o_data(mult_result_r[139][3]), .i_clk(i_clk));
Sub0000000002  u_0000000460_Sub0000000002(.i_data_1(B[139][3]), .i_data_2(C[139][3]), .o_data(mult_result_i[139][3]), .i_clk(i_clk));
Sub0000000002  u_0000000461_Sub0000000002(.i_data_1(A[140][0]), .i_data_2(B[140][0]), .o_data(mult_result_r[140][0]), .i_clk(i_clk));
Sub0000000002  u_0000000462_Sub0000000002(.i_data_1(B[140][0]), .i_data_2(C[140][0]), .o_data(mult_result_i[140][0]), .i_clk(i_clk));
Sub0000000002  u_0000000463_Sub0000000002(.i_data_1(A[140][1]), .i_data_2(B[140][1]), .o_data(mult_result_r[140][1]), .i_clk(i_clk));
Sub0000000002  u_0000000464_Sub0000000002(.i_data_1(B[140][1]), .i_data_2(C[140][1]), .o_data(mult_result_i[140][1]), .i_clk(i_clk));
Sub0000000002  u_0000000465_Sub0000000002(.i_data_1(A[140][2]), .i_data_2(B[140][2]), .o_data(mult_result_r[140][2]), .i_clk(i_clk));
Sub0000000002  u_0000000466_Sub0000000002(.i_data_1(B[140][2]), .i_data_2(C[140][2]), .o_data(mult_result_i[140][2]), .i_clk(i_clk));
Sub0000000002  u_0000000467_Sub0000000002(.i_data_1(A[140][3]), .i_data_2(B[140][3]), .o_data(mult_result_r[140][3]), .i_clk(i_clk));
Sub0000000002  u_0000000468_Sub0000000002(.i_data_1(B[140][3]), .i_data_2(C[140][3]), .o_data(mult_result_i[140][3]), .i_clk(i_clk));
Sub0000000002  u_0000000469_Sub0000000002(.i_data_1(A[141][0]), .i_data_2(B[141][0]), .o_data(mult_result_r[141][0]), .i_clk(i_clk));
Sub0000000002  u_000000046A_Sub0000000002(.i_data_1(B[141][0]), .i_data_2(C[141][0]), .o_data(mult_result_i[141][0]), .i_clk(i_clk));
Sub0000000002  u_000000046B_Sub0000000002(.i_data_1(A[141][1]), .i_data_2(B[141][1]), .o_data(mult_result_r[141][1]), .i_clk(i_clk));
Sub0000000002  u_000000046C_Sub0000000002(.i_data_1(B[141][1]), .i_data_2(C[141][1]), .o_data(mult_result_i[141][1]), .i_clk(i_clk));
Sub0000000002  u_000000046D_Sub0000000002(.i_data_1(A[141][2]), .i_data_2(B[141][2]), .o_data(mult_result_r[141][2]), .i_clk(i_clk));
Sub0000000002  u_000000046E_Sub0000000002(.i_data_1(B[141][2]), .i_data_2(C[141][2]), .o_data(mult_result_i[141][2]), .i_clk(i_clk));
Sub0000000002  u_000000046F_Sub0000000002(.i_data_1(A[141][3]), .i_data_2(B[141][3]), .o_data(mult_result_r[141][3]), .i_clk(i_clk));
Sub0000000002  u_0000000470_Sub0000000002(.i_data_1(B[141][3]), .i_data_2(C[141][3]), .o_data(mult_result_i[141][3]), .i_clk(i_clk));
Sub0000000002  u_0000000471_Sub0000000002(.i_data_1(A[142][0]), .i_data_2(B[142][0]), .o_data(mult_result_r[142][0]), .i_clk(i_clk));
Sub0000000002  u_0000000472_Sub0000000002(.i_data_1(B[142][0]), .i_data_2(C[142][0]), .o_data(mult_result_i[142][0]), .i_clk(i_clk));
Sub0000000002  u_0000000473_Sub0000000002(.i_data_1(A[142][1]), .i_data_2(B[142][1]), .o_data(mult_result_r[142][1]), .i_clk(i_clk));
Sub0000000002  u_0000000474_Sub0000000002(.i_data_1(B[142][1]), .i_data_2(C[142][1]), .o_data(mult_result_i[142][1]), .i_clk(i_clk));
Sub0000000002  u_0000000475_Sub0000000002(.i_data_1(A[142][2]), .i_data_2(B[142][2]), .o_data(mult_result_r[142][2]), .i_clk(i_clk));
Sub0000000002  u_0000000476_Sub0000000002(.i_data_1(B[142][2]), .i_data_2(C[142][2]), .o_data(mult_result_i[142][2]), .i_clk(i_clk));
Sub0000000002  u_0000000477_Sub0000000002(.i_data_1(A[142][3]), .i_data_2(B[142][3]), .o_data(mult_result_r[142][3]), .i_clk(i_clk));
Sub0000000002  u_0000000478_Sub0000000002(.i_data_1(B[142][3]), .i_data_2(C[142][3]), .o_data(mult_result_i[142][3]), .i_clk(i_clk));
Sub0000000002  u_0000000479_Sub0000000002(.i_data_1(A[143][0]), .i_data_2(B[143][0]), .o_data(mult_result_r[143][0]), .i_clk(i_clk));
Sub0000000002  u_000000047A_Sub0000000002(.i_data_1(B[143][0]), .i_data_2(C[143][0]), .o_data(mult_result_i[143][0]), .i_clk(i_clk));
Sub0000000002  u_000000047B_Sub0000000002(.i_data_1(A[143][1]), .i_data_2(B[143][1]), .o_data(mult_result_r[143][1]), .i_clk(i_clk));
Sub0000000002  u_000000047C_Sub0000000002(.i_data_1(B[143][1]), .i_data_2(C[143][1]), .o_data(mult_result_i[143][1]), .i_clk(i_clk));
Sub0000000002  u_000000047D_Sub0000000002(.i_data_1(A[143][2]), .i_data_2(B[143][2]), .o_data(mult_result_r[143][2]), .i_clk(i_clk));
Sub0000000002  u_000000047E_Sub0000000002(.i_data_1(B[143][2]), .i_data_2(C[143][2]), .o_data(mult_result_i[143][2]), .i_clk(i_clk));
Sub0000000002  u_000000047F_Sub0000000002(.i_data_1(A[143][3]), .i_data_2(B[143][3]), .o_data(mult_result_r[143][3]), .i_clk(i_clk));
Sub0000000002  u_0000000480_Sub0000000002(.i_data_1(B[143][3]), .i_data_2(C[143][3]), .o_data(mult_result_i[143][3]), .i_clk(i_clk));
Sub0000000002  u_0000000481_Sub0000000002(.i_data_1(A[144][0]), .i_data_2(B[144][0]), .o_data(mult_result_r[144][0]), .i_clk(i_clk));
Sub0000000002  u_0000000482_Sub0000000002(.i_data_1(B[144][0]), .i_data_2(C[144][0]), .o_data(mult_result_i[144][0]), .i_clk(i_clk));
Sub0000000002  u_0000000483_Sub0000000002(.i_data_1(A[144][1]), .i_data_2(B[144][1]), .o_data(mult_result_r[144][1]), .i_clk(i_clk));
Sub0000000002  u_0000000484_Sub0000000002(.i_data_1(B[144][1]), .i_data_2(C[144][1]), .o_data(mult_result_i[144][1]), .i_clk(i_clk));
Sub0000000002  u_0000000485_Sub0000000002(.i_data_1(A[144][2]), .i_data_2(B[144][2]), .o_data(mult_result_r[144][2]), .i_clk(i_clk));
Sub0000000002  u_0000000486_Sub0000000002(.i_data_1(B[144][2]), .i_data_2(C[144][2]), .o_data(mult_result_i[144][2]), .i_clk(i_clk));
Sub0000000002  u_0000000487_Sub0000000002(.i_data_1(A[144][3]), .i_data_2(B[144][3]), .o_data(mult_result_r[144][3]), .i_clk(i_clk));
Sub0000000002  u_0000000488_Sub0000000002(.i_data_1(B[144][3]), .i_data_2(C[144][3]), .o_data(mult_result_i[144][3]), .i_clk(i_clk));
Sub0000000002  u_0000000489_Sub0000000002(.i_data_1(A[145][0]), .i_data_2(B[145][0]), .o_data(mult_result_r[145][0]), .i_clk(i_clk));
Sub0000000002  u_000000048A_Sub0000000002(.i_data_1(B[145][0]), .i_data_2(C[145][0]), .o_data(mult_result_i[145][0]), .i_clk(i_clk));
Sub0000000002  u_000000048B_Sub0000000002(.i_data_1(A[145][1]), .i_data_2(B[145][1]), .o_data(mult_result_r[145][1]), .i_clk(i_clk));
Sub0000000002  u_000000048C_Sub0000000002(.i_data_1(B[145][1]), .i_data_2(C[145][1]), .o_data(mult_result_i[145][1]), .i_clk(i_clk));
Sub0000000002  u_000000048D_Sub0000000002(.i_data_1(A[145][2]), .i_data_2(B[145][2]), .o_data(mult_result_r[145][2]), .i_clk(i_clk));
Sub0000000002  u_000000048E_Sub0000000002(.i_data_1(B[145][2]), .i_data_2(C[145][2]), .o_data(mult_result_i[145][2]), .i_clk(i_clk));
Sub0000000002  u_000000048F_Sub0000000002(.i_data_1(A[145][3]), .i_data_2(B[145][3]), .o_data(mult_result_r[145][3]), .i_clk(i_clk));
Sub0000000002  u_0000000490_Sub0000000002(.i_data_1(B[145][3]), .i_data_2(C[145][3]), .o_data(mult_result_i[145][3]), .i_clk(i_clk));
Sub0000000002  u_0000000491_Sub0000000002(.i_data_1(A[146][0]), .i_data_2(B[146][0]), .o_data(mult_result_r[146][0]), .i_clk(i_clk));
Sub0000000002  u_0000000492_Sub0000000002(.i_data_1(B[146][0]), .i_data_2(C[146][0]), .o_data(mult_result_i[146][0]), .i_clk(i_clk));
Sub0000000002  u_0000000493_Sub0000000002(.i_data_1(A[146][1]), .i_data_2(B[146][1]), .o_data(mult_result_r[146][1]), .i_clk(i_clk));
Sub0000000002  u_0000000494_Sub0000000002(.i_data_1(B[146][1]), .i_data_2(C[146][1]), .o_data(mult_result_i[146][1]), .i_clk(i_clk));
Sub0000000002  u_0000000495_Sub0000000002(.i_data_1(A[146][2]), .i_data_2(B[146][2]), .o_data(mult_result_r[146][2]), .i_clk(i_clk));
Sub0000000002  u_0000000496_Sub0000000002(.i_data_1(B[146][2]), .i_data_2(C[146][2]), .o_data(mult_result_i[146][2]), .i_clk(i_clk));
Sub0000000002  u_0000000497_Sub0000000002(.i_data_1(A[146][3]), .i_data_2(B[146][3]), .o_data(mult_result_r[146][3]), .i_clk(i_clk));
Sub0000000002  u_0000000498_Sub0000000002(.i_data_1(B[146][3]), .i_data_2(C[146][3]), .o_data(mult_result_i[146][3]), .i_clk(i_clk));
Sub0000000002  u_0000000499_Sub0000000002(.i_data_1(A[147][0]), .i_data_2(B[147][0]), .o_data(mult_result_r[147][0]), .i_clk(i_clk));
Sub0000000002  u_000000049A_Sub0000000002(.i_data_1(B[147][0]), .i_data_2(C[147][0]), .o_data(mult_result_i[147][0]), .i_clk(i_clk));
Sub0000000002  u_000000049B_Sub0000000002(.i_data_1(A[147][1]), .i_data_2(B[147][1]), .o_data(mult_result_r[147][1]), .i_clk(i_clk));
Sub0000000002  u_000000049C_Sub0000000002(.i_data_1(B[147][1]), .i_data_2(C[147][1]), .o_data(mult_result_i[147][1]), .i_clk(i_clk));
Sub0000000002  u_000000049D_Sub0000000002(.i_data_1(A[147][2]), .i_data_2(B[147][2]), .o_data(mult_result_r[147][2]), .i_clk(i_clk));
Sub0000000002  u_000000049E_Sub0000000002(.i_data_1(B[147][2]), .i_data_2(C[147][2]), .o_data(mult_result_i[147][2]), .i_clk(i_clk));
Sub0000000002  u_000000049F_Sub0000000002(.i_data_1(A[147][3]), .i_data_2(B[147][3]), .o_data(mult_result_r[147][3]), .i_clk(i_clk));
Sub0000000002  u_00000004A0_Sub0000000002(.i_data_1(B[147][3]), .i_data_2(C[147][3]), .o_data(mult_result_i[147][3]), .i_clk(i_clk));
Sub0000000002  u_00000004A1_Sub0000000002(.i_data_1(A[148][0]), .i_data_2(B[148][0]), .o_data(mult_result_r[148][0]), .i_clk(i_clk));
Sub0000000002  u_00000004A2_Sub0000000002(.i_data_1(B[148][0]), .i_data_2(C[148][0]), .o_data(mult_result_i[148][0]), .i_clk(i_clk));
Sub0000000002  u_00000004A3_Sub0000000002(.i_data_1(A[148][1]), .i_data_2(B[148][1]), .o_data(mult_result_r[148][1]), .i_clk(i_clk));
Sub0000000002  u_00000004A4_Sub0000000002(.i_data_1(B[148][1]), .i_data_2(C[148][1]), .o_data(mult_result_i[148][1]), .i_clk(i_clk));
Sub0000000002  u_00000004A5_Sub0000000002(.i_data_1(A[148][2]), .i_data_2(B[148][2]), .o_data(mult_result_r[148][2]), .i_clk(i_clk));
Sub0000000002  u_00000004A6_Sub0000000002(.i_data_1(B[148][2]), .i_data_2(C[148][2]), .o_data(mult_result_i[148][2]), .i_clk(i_clk));
Sub0000000002  u_00000004A7_Sub0000000002(.i_data_1(A[148][3]), .i_data_2(B[148][3]), .o_data(mult_result_r[148][3]), .i_clk(i_clk));
Sub0000000002  u_00000004A8_Sub0000000002(.i_data_1(B[148][3]), .i_data_2(C[148][3]), .o_data(mult_result_i[148][3]), .i_clk(i_clk));
Sub0000000002  u_00000004A9_Sub0000000002(.i_data_1(A[149][0]), .i_data_2(B[149][0]), .o_data(mult_result_r[149][0]), .i_clk(i_clk));
Sub0000000002  u_00000004AA_Sub0000000002(.i_data_1(B[149][0]), .i_data_2(C[149][0]), .o_data(mult_result_i[149][0]), .i_clk(i_clk));
Sub0000000002  u_00000004AB_Sub0000000002(.i_data_1(A[149][1]), .i_data_2(B[149][1]), .o_data(mult_result_r[149][1]), .i_clk(i_clk));
Sub0000000002  u_00000004AC_Sub0000000002(.i_data_1(B[149][1]), .i_data_2(C[149][1]), .o_data(mult_result_i[149][1]), .i_clk(i_clk));
Sub0000000002  u_00000004AD_Sub0000000002(.i_data_1(A[149][2]), .i_data_2(B[149][2]), .o_data(mult_result_r[149][2]), .i_clk(i_clk));
Sub0000000002  u_00000004AE_Sub0000000002(.i_data_1(B[149][2]), .i_data_2(C[149][2]), .o_data(mult_result_i[149][2]), .i_clk(i_clk));
Sub0000000002  u_00000004AF_Sub0000000002(.i_data_1(A[149][3]), .i_data_2(B[149][3]), .o_data(mult_result_r[149][3]), .i_clk(i_clk));
Sub0000000002  u_00000004B0_Sub0000000002(.i_data_1(B[149][3]), .i_data_2(C[149][3]), .o_data(mult_result_i[149][3]), .i_clk(i_clk));
Sub0000000002  u_00000004B1_Sub0000000002(.i_data_1(A[150][0]), .i_data_2(B[150][0]), .o_data(mult_result_r[150][0]), .i_clk(i_clk));
Sub0000000002  u_00000004B2_Sub0000000002(.i_data_1(B[150][0]), .i_data_2(C[150][0]), .o_data(mult_result_i[150][0]), .i_clk(i_clk));
Sub0000000002  u_00000004B3_Sub0000000002(.i_data_1(A[150][1]), .i_data_2(B[150][1]), .o_data(mult_result_r[150][1]), .i_clk(i_clk));
Sub0000000002  u_00000004B4_Sub0000000002(.i_data_1(B[150][1]), .i_data_2(C[150][1]), .o_data(mult_result_i[150][1]), .i_clk(i_clk));
Sub0000000002  u_00000004B5_Sub0000000002(.i_data_1(A[150][2]), .i_data_2(B[150][2]), .o_data(mult_result_r[150][2]), .i_clk(i_clk));
Sub0000000002  u_00000004B6_Sub0000000002(.i_data_1(B[150][2]), .i_data_2(C[150][2]), .o_data(mult_result_i[150][2]), .i_clk(i_clk));
Sub0000000002  u_00000004B7_Sub0000000002(.i_data_1(A[150][3]), .i_data_2(B[150][3]), .o_data(mult_result_r[150][3]), .i_clk(i_clk));
Sub0000000002  u_00000004B8_Sub0000000002(.i_data_1(B[150][3]), .i_data_2(C[150][3]), .o_data(mult_result_i[150][3]), .i_clk(i_clk));
Sub0000000002  u_00000004B9_Sub0000000002(.i_data_1(A[151][0]), .i_data_2(B[151][0]), .o_data(mult_result_r[151][0]), .i_clk(i_clk));
Sub0000000002  u_00000004BA_Sub0000000002(.i_data_1(B[151][0]), .i_data_2(C[151][0]), .o_data(mult_result_i[151][0]), .i_clk(i_clk));
Sub0000000002  u_00000004BB_Sub0000000002(.i_data_1(A[151][1]), .i_data_2(B[151][1]), .o_data(mult_result_r[151][1]), .i_clk(i_clk));
Sub0000000002  u_00000004BC_Sub0000000002(.i_data_1(B[151][1]), .i_data_2(C[151][1]), .o_data(mult_result_i[151][1]), .i_clk(i_clk));
Sub0000000002  u_00000004BD_Sub0000000002(.i_data_1(A[151][2]), .i_data_2(B[151][2]), .o_data(mult_result_r[151][2]), .i_clk(i_clk));
Sub0000000002  u_00000004BE_Sub0000000002(.i_data_1(B[151][2]), .i_data_2(C[151][2]), .o_data(mult_result_i[151][2]), .i_clk(i_clk));
Sub0000000002  u_00000004BF_Sub0000000002(.i_data_1(A[151][3]), .i_data_2(B[151][3]), .o_data(mult_result_r[151][3]), .i_clk(i_clk));
Sub0000000002  u_00000004C0_Sub0000000002(.i_data_1(B[151][3]), .i_data_2(C[151][3]), .o_data(mult_result_i[151][3]), .i_clk(i_clk));
Sub0000000002  u_00000004C1_Sub0000000002(.i_data_1(A[152][0]), .i_data_2(B[152][0]), .o_data(mult_result_r[152][0]), .i_clk(i_clk));
Sub0000000002  u_00000004C2_Sub0000000002(.i_data_1(B[152][0]), .i_data_2(C[152][0]), .o_data(mult_result_i[152][0]), .i_clk(i_clk));
Sub0000000002  u_00000004C3_Sub0000000002(.i_data_1(A[152][1]), .i_data_2(B[152][1]), .o_data(mult_result_r[152][1]), .i_clk(i_clk));
Sub0000000002  u_00000004C4_Sub0000000002(.i_data_1(B[152][1]), .i_data_2(C[152][1]), .o_data(mult_result_i[152][1]), .i_clk(i_clk));
Sub0000000002  u_00000004C5_Sub0000000002(.i_data_1(A[152][2]), .i_data_2(B[152][2]), .o_data(mult_result_r[152][2]), .i_clk(i_clk));
Sub0000000002  u_00000004C6_Sub0000000002(.i_data_1(B[152][2]), .i_data_2(C[152][2]), .o_data(mult_result_i[152][2]), .i_clk(i_clk));
Sub0000000002  u_00000004C7_Sub0000000002(.i_data_1(A[152][3]), .i_data_2(B[152][3]), .o_data(mult_result_r[152][3]), .i_clk(i_clk));
Sub0000000002  u_00000004C8_Sub0000000002(.i_data_1(B[152][3]), .i_data_2(C[152][3]), .o_data(mult_result_i[152][3]), .i_clk(i_clk));
Sub0000000002  u_00000004C9_Sub0000000002(.i_data_1(A[153][0]), .i_data_2(B[153][0]), .o_data(mult_result_r[153][0]), .i_clk(i_clk));
Sub0000000002  u_00000004CA_Sub0000000002(.i_data_1(B[153][0]), .i_data_2(C[153][0]), .o_data(mult_result_i[153][0]), .i_clk(i_clk));
Sub0000000002  u_00000004CB_Sub0000000002(.i_data_1(A[153][1]), .i_data_2(B[153][1]), .o_data(mult_result_r[153][1]), .i_clk(i_clk));
Sub0000000002  u_00000004CC_Sub0000000002(.i_data_1(B[153][1]), .i_data_2(C[153][1]), .o_data(mult_result_i[153][1]), .i_clk(i_clk));
Sub0000000002  u_00000004CD_Sub0000000002(.i_data_1(A[153][2]), .i_data_2(B[153][2]), .o_data(mult_result_r[153][2]), .i_clk(i_clk));
Sub0000000002  u_00000004CE_Sub0000000002(.i_data_1(B[153][2]), .i_data_2(C[153][2]), .o_data(mult_result_i[153][2]), .i_clk(i_clk));
Sub0000000002  u_00000004CF_Sub0000000002(.i_data_1(A[153][3]), .i_data_2(B[153][3]), .o_data(mult_result_r[153][3]), .i_clk(i_clk));
Sub0000000002  u_00000004D0_Sub0000000002(.i_data_1(B[153][3]), .i_data_2(C[153][3]), .o_data(mult_result_i[153][3]), .i_clk(i_clk));
Sub0000000002  u_00000004D1_Sub0000000002(.i_data_1(A[154][0]), .i_data_2(B[154][0]), .o_data(mult_result_r[154][0]), .i_clk(i_clk));
Sub0000000002  u_00000004D2_Sub0000000002(.i_data_1(B[154][0]), .i_data_2(C[154][0]), .o_data(mult_result_i[154][0]), .i_clk(i_clk));
Sub0000000002  u_00000004D3_Sub0000000002(.i_data_1(A[154][1]), .i_data_2(B[154][1]), .o_data(mult_result_r[154][1]), .i_clk(i_clk));
Sub0000000002  u_00000004D4_Sub0000000002(.i_data_1(B[154][1]), .i_data_2(C[154][1]), .o_data(mult_result_i[154][1]), .i_clk(i_clk));
Sub0000000002  u_00000004D5_Sub0000000002(.i_data_1(A[154][2]), .i_data_2(B[154][2]), .o_data(mult_result_r[154][2]), .i_clk(i_clk));
Sub0000000002  u_00000004D6_Sub0000000002(.i_data_1(B[154][2]), .i_data_2(C[154][2]), .o_data(mult_result_i[154][2]), .i_clk(i_clk));
Sub0000000002  u_00000004D7_Sub0000000002(.i_data_1(A[154][3]), .i_data_2(B[154][3]), .o_data(mult_result_r[154][3]), .i_clk(i_clk));
Sub0000000002  u_00000004D8_Sub0000000002(.i_data_1(B[154][3]), .i_data_2(C[154][3]), .o_data(mult_result_i[154][3]), .i_clk(i_clk));
Sub0000000002  u_00000004D9_Sub0000000002(.i_data_1(A[155][0]), .i_data_2(B[155][0]), .o_data(mult_result_r[155][0]), .i_clk(i_clk));
Sub0000000002  u_00000004DA_Sub0000000002(.i_data_1(B[155][0]), .i_data_2(C[155][0]), .o_data(mult_result_i[155][0]), .i_clk(i_clk));
Sub0000000002  u_00000004DB_Sub0000000002(.i_data_1(A[155][1]), .i_data_2(B[155][1]), .o_data(mult_result_r[155][1]), .i_clk(i_clk));
Sub0000000002  u_00000004DC_Sub0000000002(.i_data_1(B[155][1]), .i_data_2(C[155][1]), .o_data(mult_result_i[155][1]), .i_clk(i_clk));
Sub0000000002  u_00000004DD_Sub0000000002(.i_data_1(A[155][2]), .i_data_2(B[155][2]), .o_data(mult_result_r[155][2]), .i_clk(i_clk));
Sub0000000002  u_00000004DE_Sub0000000002(.i_data_1(B[155][2]), .i_data_2(C[155][2]), .o_data(mult_result_i[155][2]), .i_clk(i_clk));
Sub0000000002  u_00000004DF_Sub0000000002(.i_data_1(A[155][3]), .i_data_2(B[155][3]), .o_data(mult_result_r[155][3]), .i_clk(i_clk));
Sub0000000002  u_00000004E0_Sub0000000002(.i_data_1(B[155][3]), .i_data_2(C[155][3]), .o_data(mult_result_i[155][3]), .i_clk(i_clk));
Sub0000000002  u_00000004E1_Sub0000000002(.i_data_1(A[156][0]), .i_data_2(B[156][0]), .o_data(mult_result_r[156][0]), .i_clk(i_clk));
Sub0000000002  u_00000004E2_Sub0000000002(.i_data_1(B[156][0]), .i_data_2(C[156][0]), .o_data(mult_result_i[156][0]), .i_clk(i_clk));
Sub0000000002  u_00000004E3_Sub0000000002(.i_data_1(A[156][1]), .i_data_2(B[156][1]), .o_data(mult_result_r[156][1]), .i_clk(i_clk));
Sub0000000002  u_00000004E4_Sub0000000002(.i_data_1(B[156][1]), .i_data_2(C[156][1]), .o_data(mult_result_i[156][1]), .i_clk(i_clk));
Sub0000000002  u_00000004E5_Sub0000000002(.i_data_1(A[156][2]), .i_data_2(B[156][2]), .o_data(mult_result_r[156][2]), .i_clk(i_clk));
Sub0000000002  u_00000004E6_Sub0000000002(.i_data_1(B[156][2]), .i_data_2(C[156][2]), .o_data(mult_result_i[156][2]), .i_clk(i_clk));
Sub0000000002  u_00000004E7_Sub0000000002(.i_data_1(A[156][3]), .i_data_2(B[156][3]), .o_data(mult_result_r[156][3]), .i_clk(i_clk));
Sub0000000002  u_00000004E8_Sub0000000002(.i_data_1(B[156][3]), .i_data_2(C[156][3]), .o_data(mult_result_i[156][3]), .i_clk(i_clk));
Sub0000000002  u_00000004E9_Sub0000000002(.i_data_1(A[157][0]), .i_data_2(B[157][0]), .o_data(mult_result_r[157][0]), .i_clk(i_clk));
Sub0000000002  u_00000004EA_Sub0000000002(.i_data_1(B[157][0]), .i_data_2(C[157][0]), .o_data(mult_result_i[157][0]), .i_clk(i_clk));
Sub0000000002  u_00000004EB_Sub0000000002(.i_data_1(A[157][1]), .i_data_2(B[157][1]), .o_data(mult_result_r[157][1]), .i_clk(i_clk));
Sub0000000002  u_00000004EC_Sub0000000002(.i_data_1(B[157][1]), .i_data_2(C[157][1]), .o_data(mult_result_i[157][1]), .i_clk(i_clk));
Sub0000000002  u_00000004ED_Sub0000000002(.i_data_1(A[157][2]), .i_data_2(B[157][2]), .o_data(mult_result_r[157][2]), .i_clk(i_clk));
Sub0000000002  u_00000004EE_Sub0000000002(.i_data_1(B[157][2]), .i_data_2(C[157][2]), .o_data(mult_result_i[157][2]), .i_clk(i_clk));
Sub0000000002  u_00000004EF_Sub0000000002(.i_data_1(A[157][3]), .i_data_2(B[157][3]), .o_data(mult_result_r[157][3]), .i_clk(i_clk));
Sub0000000002  u_00000004F0_Sub0000000002(.i_data_1(B[157][3]), .i_data_2(C[157][3]), .o_data(mult_result_i[157][3]), .i_clk(i_clk));
Sub0000000002  u_00000004F1_Sub0000000002(.i_data_1(A[158][0]), .i_data_2(B[158][0]), .o_data(mult_result_r[158][0]), .i_clk(i_clk));
Sub0000000002  u_00000004F2_Sub0000000002(.i_data_1(B[158][0]), .i_data_2(C[158][0]), .o_data(mult_result_i[158][0]), .i_clk(i_clk));
Sub0000000002  u_00000004F3_Sub0000000002(.i_data_1(A[158][1]), .i_data_2(B[158][1]), .o_data(mult_result_r[158][1]), .i_clk(i_clk));
Sub0000000002  u_00000004F4_Sub0000000002(.i_data_1(B[158][1]), .i_data_2(C[158][1]), .o_data(mult_result_i[158][1]), .i_clk(i_clk));
Sub0000000002  u_00000004F5_Sub0000000002(.i_data_1(A[158][2]), .i_data_2(B[158][2]), .o_data(mult_result_r[158][2]), .i_clk(i_clk));
Sub0000000002  u_00000004F6_Sub0000000002(.i_data_1(B[158][2]), .i_data_2(C[158][2]), .o_data(mult_result_i[158][2]), .i_clk(i_clk));
Sub0000000002  u_00000004F7_Sub0000000002(.i_data_1(A[158][3]), .i_data_2(B[158][3]), .o_data(mult_result_r[158][3]), .i_clk(i_clk));
Sub0000000002  u_00000004F8_Sub0000000002(.i_data_1(B[158][3]), .i_data_2(C[158][3]), .o_data(mult_result_i[158][3]), .i_clk(i_clk));
Sub0000000002  u_00000004F9_Sub0000000002(.i_data_1(A[159][0]), .i_data_2(B[159][0]), .o_data(mult_result_r[159][0]), .i_clk(i_clk));
Sub0000000002  u_00000004FA_Sub0000000002(.i_data_1(B[159][0]), .i_data_2(C[159][0]), .o_data(mult_result_i[159][0]), .i_clk(i_clk));
Sub0000000002  u_00000004FB_Sub0000000002(.i_data_1(A[159][1]), .i_data_2(B[159][1]), .o_data(mult_result_r[159][1]), .i_clk(i_clk));
Sub0000000002  u_00000004FC_Sub0000000002(.i_data_1(B[159][1]), .i_data_2(C[159][1]), .o_data(mult_result_i[159][1]), .i_clk(i_clk));
Sub0000000002  u_00000004FD_Sub0000000002(.i_data_1(A[159][2]), .i_data_2(B[159][2]), .o_data(mult_result_r[159][2]), .i_clk(i_clk));
Sub0000000002  u_00000004FE_Sub0000000002(.i_data_1(B[159][2]), .i_data_2(C[159][2]), .o_data(mult_result_i[159][2]), .i_clk(i_clk));
Sub0000000002  u_00000004FF_Sub0000000002(.i_data_1(A[159][3]), .i_data_2(B[159][3]), .o_data(mult_result_r[159][3]), .i_clk(i_clk));
Sub0000000002  u_0000000500_Sub0000000002(.i_data_1(B[159][3]), .i_data_2(C[159][3]), .o_data(mult_result_i[159][3]), .i_clk(i_clk));
Sub0000000002  u_0000000501_Sub0000000002(.i_data_1(A[160][0]), .i_data_2(B[160][0]), .o_data(mult_result_r[160][0]), .i_clk(i_clk));
Sub0000000002  u_0000000502_Sub0000000002(.i_data_1(B[160][0]), .i_data_2(C[160][0]), .o_data(mult_result_i[160][0]), .i_clk(i_clk));
Sub0000000002  u_0000000503_Sub0000000002(.i_data_1(A[160][1]), .i_data_2(B[160][1]), .o_data(mult_result_r[160][1]), .i_clk(i_clk));
Sub0000000002  u_0000000504_Sub0000000002(.i_data_1(B[160][1]), .i_data_2(C[160][1]), .o_data(mult_result_i[160][1]), .i_clk(i_clk));
Sub0000000002  u_0000000505_Sub0000000002(.i_data_1(A[160][2]), .i_data_2(B[160][2]), .o_data(mult_result_r[160][2]), .i_clk(i_clk));
Sub0000000002  u_0000000506_Sub0000000002(.i_data_1(B[160][2]), .i_data_2(C[160][2]), .o_data(mult_result_i[160][2]), .i_clk(i_clk));
Sub0000000002  u_0000000507_Sub0000000002(.i_data_1(A[160][3]), .i_data_2(B[160][3]), .o_data(mult_result_r[160][3]), .i_clk(i_clk));
Sub0000000002  u_0000000508_Sub0000000002(.i_data_1(B[160][3]), .i_data_2(C[160][3]), .o_data(mult_result_i[160][3]), .i_clk(i_clk));
Sub0000000002  u_0000000509_Sub0000000002(.i_data_1(A[161][0]), .i_data_2(B[161][0]), .o_data(mult_result_r[161][0]), .i_clk(i_clk));
Sub0000000002  u_000000050A_Sub0000000002(.i_data_1(B[161][0]), .i_data_2(C[161][0]), .o_data(mult_result_i[161][0]), .i_clk(i_clk));
Sub0000000002  u_000000050B_Sub0000000002(.i_data_1(A[161][1]), .i_data_2(B[161][1]), .o_data(mult_result_r[161][1]), .i_clk(i_clk));
Sub0000000002  u_000000050C_Sub0000000002(.i_data_1(B[161][1]), .i_data_2(C[161][1]), .o_data(mult_result_i[161][1]), .i_clk(i_clk));
Sub0000000002  u_000000050D_Sub0000000002(.i_data_1(A[161][2]), .i_data_2(B[161][2]), .o_data(mult_result_r[161][2]), .i_clk(i_clk));
Sub0000000002  u_000000050E_Sub0000000002(.i_data_1(B[161][2]), .i_data_2(C[161][2]), .o_data(mult_result_i[161][2]), .i_clk(i_clk));
Sub0000000002  u_000000050F_Sub0000000002(.i_data_1(A[161][3]), .i_data_2(B[161][3]), .o_data(mult_result_r[161][3]), .i_clk(i_clk));
Sub0000000002  u_0000000510_Sub0000000002(.i_data_1(B[161][3]), .i_data_2(C[161][3]), .o_data(mult_result_i[161][3]), .i_clk(i_clk));
Sub0000000002  u_0000000511_Sub0000000002(.i_data_1(A[162][0]), .i_data_2(B[162][0]), .o_data(mult_result_r[162][0]), .i_clk(i_clk));
Sub0000000002  u_0000000512_Sub0000000002(.i_data_1(B[162][0]), .i_data_2(C[162][0]), .o_data(mult_result_i[162][0]), .i_clk(i_clk));
Sub0000000002  u_0000000513_Sub0000000002(.i_data_1(A[162][1]), .i_data_2(B[162][1]), .o_data(mult_result_r[162][1]), .i_clk(i_clk));
Sub0000000002  u_0000000514_Sub0000000002(.i_data_1(B[162][1]), .i_data_2(C[162][1]), .o_data(mult_result_i[162][1]), .i_clk(i_clk));
Sub0000000002  u_0000000515_Sub0000000002(.i_data_1(A[162][2]), .i_data_2(B[162][2]), .o_data(mult_result_r[162][2]), .i_clk(i_clk));
Sub0000000002  u_0000000516_Sub0000000002(.i_data_1(B[162][2]), .i_data_2(C[162][2]), .o_data(mult_result_i[162][2]), .i_clk(i_clk));
Sub0000000002  u_0000000517_Sub0000000002(.i_data_1(A[162][3]), .i_data_2(B[162][3]), .o_data(mult_result_r[162][3]), .i_clk(i_clk));
Sub0000000002  u_0000000518_Sub0000000002(.i_data_1(B[162][3]), .i_data_2(C[162][3]), .o_data(mult_result_i[162][3]), .i_clk(i_clk));
Sub0000000002  u_0000000519_Sub0000000002(.i_data_1(A[163][0]), .i_data_2(B[163][0]), .o_data(mult_result_r[163][0]), .i_clk(i_clk));
Sub0000000002  u_000000051A_Sub0000000002(.i_data_1(B[163][0]), .i_data_2(C[163][0]), .o_data(mult_result_i[163][0]), .i_clk(i_clk));
Sub0000000002  u_000000051B_Sub0000000002(.i_data_1(A[163][1]), .i_data_2(B[163][1]), .o_data(mult_result_r[163][1]), .i_clk(i_clk));
Sub0000000002  u_000000051C_Sub0000000002(.i_data_1(B[163][1]), .i_data_2(C[163][1]), .o_data(mult_result_i[163][1]), .i_clk(i_clk));
Sub0000000002  u_000000051D_Sub0000000002(.i_data_1(A[163][2]), .i_data_2(B[163][2]), .o_data(mult_result_r[163][2]), .i_clk(i_clk));
Sub0000000002  u_000000051E_Sub0000000002(.i_data_1(B[163][2]), .i_data_2(C[163][2]), .o_data(mult_result_i[163][2]), .i_clk(i_clk));
Sub0000000002  u_000000051F_Sub0000000002(.i_data_1(A[163][3]), .i_data_2(B[163][3]), .o_data(mult_result_r[163][3]), .i_clk(i_clk));
Sub0000000002  u_0000000520_Sub0000000002(.i_data_1(B[163][3]), .i_data_2(C[163][3]), .o_data(mult_result_i[163][3]), .i_clk(i_clk));
Sub0000000002  u_0000000521_Sub0000000002(.i_data_1(A[164][0]), .i_data_2(B[164][0]), .o_data(mult_result_r[164][0]), .i_clk(i_clk));
Sub0000000002  u_0000000522_Sub0000000002(.i_data_1(B[164][0]), .i_data_2(C[164][0]), .o_data(mult_result_i[164][0]), .i_clk(i_clk));
Sub0000000002  u_0000000523_Sub0000000002(.i_data_1(A[164][1]), .i_data_2(B[164][1]), .o_data(mult_result_r[164][1]), .i_clk(i_clk));
Sub0000000002  u_0000000524_Sub0000000002(.i_data_1(B[164][1]), .i_data_2(C[164][1]), .o_data(mult_result_i[164][1]), .i_clk(i_clk));
Sub0000000002  u_0000000525_Sub0000000002(.i_data_1(A[164][2]), .i_data_2(B[164][2]), .o_data(mult_result_r[164][2]), .i_clk(i_clk));
Sub0000000002  u_0000000526_Sub0000000002(.i_data_1(B[164][2]), .i_data_2(C[164][2]), .o_data(mult_result_i[164][2]), .i_clk(i_clk));
Sub0000000002  u_0000000527_Sub0000000002(.i_data_1(A[164][3]), .i_data_2(B[164][3]), .o_data(mult_result_r[164][3]), .i_clk(i_clk));
Sub0000000002  u_0000000528_Sub0000000002(.i_data_1(B[164][3]), .i_data_2(C[164][3]), .o_data(mult_result_i[164][3]), .i_clk(i_clk));
Sub0000000002  u_0000000529_Sub0000000002(.i_data_1(A[165][0]), .i_data_2(B[165][0]), .o_data(mult_result_r[165][0]), .i_clk(i_clk));
Sub0000000002  u_000000052A_Sub0000000002(.i_data_1(B[165][0]), .i_data_2(C[165][0]), .o_data(mult_result_i[165][0]), .i_clk(i_clk));
Sub0000000002  u_000000052B_Sub0000000002(.i_data_1(A[165][1]), .i_data_2(B[165][1]), .o_data(mult_result_r[165][1]), .i_clk(i_clk));
Sub0000000002  u_000000052C_Sub0000000002(.i_data_1(B[165][1]), .i_data_2(C[165][1]), .o_data(mult_result_i[165][1]), .i_clk(i_clk));
Sub0000000002  u_000000052D_Sub0000000002(.i_data_1(A[165][2]), .i_data_2(B[165][2]), .o_data(mult_result_r[165][2]), .i_clk(i_clk));
Sub0000000002  u_000000052E_Sub0000000002(.i_data_1(B[165][2]), .i_data_2(C[165][2]), .o_data(mult_result_i[165][2]), .i_clk(i_clk));
Sub0000000002  u_000000052F_Sub0000000002(.i_data_1(A[165][3]), .i_data_2(B[165][3]), .o_data(mult_result_r[165][3]), .i_clk(i_clk));
Sub0000000002  u_0000000530_Sub0000000002(.i_data_1(B[165][3]), .i_data_2(C[165][3]), .o_data(mult_result_i[165][3]), .i_clk(i_clk));
Sub0000000002  u_0000000531_Sub0000000002(.i_data_1(A[166][0]), .i_data_2(B[166][0]), .o_data(mult_result_r[166][0]), .i_clk(i_clk));
Sub0000000002  u_0000000532_Sub0000000002(.i_data_1(B[166][0]), .i_data_2(C[166][0]), .o_data(mult_result_i[166][0]), .i_clk(i_clk));
Sub0000000002  u_0000000533_Sub0000000002(.i_data_1(A[166][1]), .i_data_2(B[166][1]), .o_data(mult_result_r[166][1]), .i_clk(i_clk));
Sub0000000002  u_0000000534_Sub0000000002(.i_data_1(B[166][1]), .i_data_2(C[166][1]), .o_data(mult_result_i[166][1]), .i_clk(i_clk));
Sub0000000002  u_0000000535_Sub0000000002(.i_data_1(A[166][2]), .i_data_2(B[166][2]), .o_data(mult_result_r[166][2]), .i_clk(i_clk));
Sub0000000002  u_0000000536_Sub0000000002(.i_data_1(B[166][2]), .i_data_2(C[166][2]), .o_data(mult_result_i[166][2]), .i_clk(i_clk));
Sub0000000002  u_0000000537_Sub0000000002(.i_data_1(A[166][3]), .i_data_2(B[166][3]), .o_data(mult_result_r[166][3]), .i_clk(i_clk));
Sub0000000002  u_0000000538_Sub0000000002(.i_data_1(B[166][3]), .i_data_2(C[166][3]), .o_data(mult_result_i[166][3]), .i_clk(i_clk));
Sub0000000002  u_0000000539_Sub0000000002(.i_data_1(A[167][0]), .i_data_2(B[167][0]), .o_data(mult_result_r[167][0]), .i_clk(i_clk));
Sub0000000002  u_000000053A_Sub0000000002(.i_data_1(B[167][0]), .i_data_2(C[167][0]), .o_data(mult_result_i[167][0]), .i_clk(i_clk));
Sub0000000002  u_000000053B_Sub0000000002(.i_data_1(A[167][1]), .i_data_2(B[167][1]), .o_data(mult_result_r[167][1]), .i_clk(i_clk));
Sub0000000002  u_000000053C_Sub0000000002(.i_data_1(B[167][1]), .i_data_2(C[167][1]), .o_data(mult_result_i[167][1]), .i_clk(i_clk));
Sub0000000002  u_000000053D_Sub0000000002(.i_data_1(A[167][2]), .i_data_2(B[167][2]), .o_data(mult_result_r[167][2]), .i_clk(i_clk));
Sub0000000002  u_000000053E_Sub0000000002(.i_data_1(B[167][2]), .i_data_2(C[167][2]), .o_data(mult_result_i[167][2]), .i_clk(i_clk));
Sub0000000002  u_000000053F_Sub0000000002(.i_data_1(A[167][3]), .i_data_2(B[167][3]), .o_data(mult_result_r[167][3]), .i_clk(i_clk));
Sub0000000002  u_0000000540_Sub0000000002(.i_data_1(B[167][3]), .i_data_2(C[167][3]), .o_data(mult_result_i[167][3]), .i_clk(i_clk));
Sub0000000002  u_0000000541_Sub0000000002(.i_data_1(A[168][0]), .i_data_2(B[168][0]), .o_data(mult_result_r[168][0]), .i_clk(i_clk));
Sub0000000002  u_0000000542_Sub0000000002(.i_data_1(B[168][0]), .i_data_2(C[168][0]), .o_data(mult_result_i[168][0]), .i_clk(i_clk));
Sub0000000002  u_0000000543_Sub0000000002(.i_data_1(A[168][1]), .i_data_2(B[168][1]), .o_data(mult_result_r[168][1]), .i_clk(i_clk));
Sub0000000002  u_0000000544_Sub0000000002(.i_data_1(B[168][1]), .i_data_2(C[168][1]), .o_data(mult_result_i[168][1]), .i_clk(i_clk));
Sub0000000002  u_0000000545_Sub0000000002(.i_data_1(A[168][2]), .i_data_2(B[168][2]), .o_data(mult_result_r[168][2]), .i_clk(i_clk));
Sub0000000002  u_0000000546_Sub0000000002(.i_data_1(B[168][2]), .i_data_2(C[168][2]), .o_data(mult_result_i[168][2]), .i_clk(i_clk));
Sub0000000002  u_0000000547_Sub0000000002(.i_data_1(A[168][3]), .i_data_2(B[168][3]), .o_data(mult_result_r[168][3]), .i_clk(i_clk));
Sub0000000002  u_0000000548_Sub0000000002(.i_data_1(B[168][3]), .i_data_2(C[168][3]), .o_data(mult_result_i[168][3]), .i_clk(i_clk));
Sub0000000002  u_0000000549_Sub0000000002(.i_data_1(A[169][0]), .i_data_2(B[169][0]), .o_data(mult_result_r[169][0]), .i_clk(i_clk));
Sub0000000002  u_000000054A_Sub0000000002(.i_data_1(B[169][0]), .i_data_2(C[169][0]), .o_data(mult_result_i[169][0]), .i_clk(i_clk));
Sub0000000002  u_000000054B_Sub0000000002(.i_data_1(A[169][1]), .i_data_2(B[169][1]), .o_data(mult_result_r[169][1]), .i_clk(i_clk));
Sub0000000002  u_000000054C_Sub0000000002(.i_data_1(B[169][1]), .i_data_2(C[169][1]), .o_data(mult_result_i[169][1]), .i_clk(i_clk));
Sub0000000002  u_000000054D_Sub0000000002(.i_data_1(A[169][2]), .i_data_2(B[169][2]), .o_data(mult_result_r[169][2]), .i_clk(i_clk));
Sub0000000002  u_000000054E_Sub0000000002(.i_data_1(B[169][2]), .i_data_2(C[169][2]), .o_data(mult_result_i[169][2]), .i_clk(i_clk));
Sub0000000002  u_000000054F_Sub0000000002(.i_data_1(A[169][3]), .i_data_2(B[169][3]), .o_data(mult_result_r[169][3]), .i_clk(i_clk));
Sub0000000002  u_0000000550_Sub0000000002(.i_data_1(B[169][3]), .i_data_2(C[169][3]), .o_data(mult_result_i[169][3]), .i_clk(i_clk));
Sub0000000002  u_0000000551_Sub0000000002(.i_data_1(A[170][0]), .i_data_2(B[170][0]), .o_data(mult_result_r[170][0]), .i_clk(i_clk));
Sub0000000002  u_0000000552_Sub0000000002(.i_data_1(B[170][0]), .i_data_2(C[170][0]), .o_data(mult_result_i[170][0]), .i_clk(i_clk));
Sub0000000002  u_0000000553_Sub0000000002(.i_data_1(A[170][1]), .i_data_2(B[170][1]), .o_data(mult_result_r[170][1]), .i_clk(i_clk));
Sub0000000002  u_0000000554_Sub0000000002(.i_data_1(B[170][1]), .i_data_2(C[170][1]), .o_data(mult_result_i[170][1]), .i_clk(i_clk));
Sub0000000002  u_0000000555_Sub0000000002(.i_data_1(A[170][2]), .i_data_2(B[170][2]), .o_data(mult_result_r[170][2]), .i_clk(i_clk));
Sub0000000002  u_0000000556_Sub0000000002(.i_data_1(B[170][2]), .i_data_2(C[170][2]), .o_data(mult_result_i[170][2]), .i_clk(i_clk));
Sub0000000002  u_0000000557_Sub0000000002(.i_data_1(A[170][3]), .i_data_2(B[170][3]), .o_data(mult_result_r[170][3]), .i_clk(i_clk));
Sub0000000002  u_0000000558_Sub0000000002(.i_data_1(B[170][3]), .i_data_2(C[170][3]), .o_data(mult_result_i[170][3]), .i_clk(i_clk));
Sub0000000002  u_0000000559_Sub0000000002(.i_data_1(A[171][0]), .i_data_2(B[171][0]), .o_data(mult_result_r[171][0]), .i_clk(i_clk));
Sub0000000002  u_000000055A_Sub0000000002(.i_data_1(B[171][0]), .i_data_2(C[171][0]), .o_data(mult_result_i[171][0]), .i_clk(i_clk));
Sub0000000002  u_000000055B_Sub0000000002(.i_data_1(A[171][1]), .i_data_2(B[171][1]), .o_data(mult_result_r[171][1]), .i_clk(i_clk));
Sub0000000002  u_000000055C_Sub0000000002(.i_data_1(B[171][1]), .i_data_2(C[171][1]), .o_data(mult_result_i[171][1]), .i_clk(i_clk));
Sub0000000002  u_000000055D_Sub0000000002(.i_data_1(A[171][2]), .i_data_2(B[171][2]), .o_data(mult_result_r[171][2]), .i_clk(i_clk));
Sub0000000002  u_000000055E_Sub0000000002(.i_data_1(B[171][2]), .i_data_2(C[171][2]), .o_data(mult_result_i[171][2]), .i_clk(i_clk));
Sub0000000002  u_000000055F_Sub0000000002(.i_data_1(A[171][3]), .i_data_2(B[171][3]), .o_data(mult_result_r[171][3]), .i_clk(i_clk));
Sub0000000002  u_0000000560_Sub0000000002(.i_data_1(B[171][3]), .i_data_2(C[171][3]), .o_data(mult_result_i[171][3]), .i_clk(i_clk));
Sub0000000002  u_0000000561_Sub0000000002(.i_data_1(A[172][0]), .i_data_2(B[172][0]), .o_data(mult_result_r[172][0]), .i_clk(i_clk));
Sub0000000002  u_0000000562_Sub0000000002(.i_data_1(B[172][0]), .i_data_2(C[172][0]), .o_data(mult_result_i[172][0]), .i_clk(i_clk));
Sub0000000002  u_0000000563_Sub0000000002(.i_data_1(A[172][1]), .i_data_2(B[172][1]), .o_data(mult_result_r[172][1]), .i_clk(i_clk));
Sub0000000002  u_0000000564_Sub0000000002(.i_data_1(B[172][1]), .i_data_2(C[172][1]), .o_data(mult_result_i[172][1]), .i_clk(i_clk));
Sub0000000002  u_0000000565_Sub0000000002(.i_data_1(A[172][2]), .i_data_2(B[172][2]), .o_data(mult_result_r[172][2]), .i_clk(i_clk));
Sub0000000002  u_0000000566_Sub0000000002(.i_data_1(B[172][2]), .i_data_2(C[172][2]), .o_data(mult_result_i[172][2]), .i_clk(i_clk));
Sub0000000002  u_0000000567_Sub0000000002(.i_data_1(A[172][3]), .i_data_2(B[172][3]), .o_data(mult_result_r[172][3]), .i_clk(i_clk));
Sub0000000002  u_0000000568_Sub0000000002(.i_data_1(B[172][3]), .i_data_2(C[172][3]), .o_data(mult_result_i[172][3]), .i_clk(i_clk));
Sub0000000002  u_0000000569_Sub0000000002(.i_data_1(A[173][0]), .i_data_2(B[173][0]), .o_data(mult_result_r[173][0]), .i_clk(i_clk));
Sub0000000002  u_000000056A_Sub0000000002(.i_data_1(B[173][0]), .i_data_2(C[173][0]), .o_data(mult_result_i[173][0]), .i_clk(i_clk));
Sub0000000002  u_000000056B_Sub0000000002(.i_data_1(A[173][1]), .i_data_2(B[173][1]), .o_data(mult_result_r[173][1]), .i_clk(i_clk));
Sub0000000002  u_000000056C_Sub0000000002(.i_data_1(B[173][1]), .i_data_2(C[173][1]), .o_data(mult_result_i[173][1]), .i_clk(i_clk));
Sub0000000002  u_000000056D_Sub0000000002(.i_data_1(A[173][2]), .i_data_2(B[173][2]), .o_data(mult_result_r[173][2]), .i_clk(i_clk));
Sub0000000002  u_000000056E_Sub0000000002(.i_data_1(B[173][2]), .i_data_2(C[173][2]), .o_data(mult_result_i[173][2]), .i_clk(i_clk));
Sub0000000002  u_000000056F_Sub0000000002(.i_data_1(A[173][3]), .i_data_2(B[173][3]), .o_data(mult_result_r[173][3]), .i_clk(i_clk));
Sub0000000002  u_0000000570_Sub0000000002(.i_data_1(B[173][3]), .i_data_2(C[173][3]), .o_data(mult_result_i[173][3]), .i_clk(i_clk));
Sub0000000002  u_0000000571_Sub0000000002(.i_data_1(A[174][0]), .i_data_2(B[174][0]), .o_data(mult_result_r[174][0]), .i_clk(i_clk));
Sub0000000002  u_0000000572_Sub0000000002(.i_data_1(B[174][0]), .i_data_2(C[174][0]), .o_data(mult_result_i[174][0]), .i_clk(i_clk));
Sub0000000002  u_0000000573_Sub0000000002(.i_data_1(A[174][1]), .i_data_2(B[174][1]), .o_data(mult_result_r[174][1]), .i_clk(i_clk));
Sub0000000002  u_0000000574_Sub0000000002(.i_data_1(B[174][1]), .i_data_2(C[174][1]), .o_data(mult_result_i[174][1]), .i_clk(i_clk));
Sub0000000002  u_0000000575_Sub0000000002(.i_data_1(A[174][2]), .i_data_2(B[174][2]), .o_data(mult_result_r[174][2]), .i_clk(i_clk));
Sub0000000002  u_0000000576_Sub0000000002(.i_data_1(B[174][2]), .i_data_2(C[174][2]), .o_data(mult_result_i[174][2]), .i_clk(i_clk));
Sub0000000002  u_0000000577_Sub0000000002(.i_data_1(A[174][3]), .i_data_2(B[174][3]), .o_data(mult_result_r[174][3]), .i_clk(i_clk));
Sub0000000002  u_0000000578_Sub0000000002(.i_data_1(B[174][3]), .i_data_2(C[174][3]), .o_data(mult_result_i[174][3]), .i_clk(i_clk));
Sub0000000002  u_0000000579_Sub0000000002(.i_data_1(A[175][0]), .i_data_2(B[175][0]), .o_data(mult_result_r[175][0]), .i_clk(i_clk));
Sub0000000002  u_000000057A_Sub0000000002(.i_data_1(B[175][0]), .i_data_2(C[175][0]), .o_data(mult_result_i[175][0]), .i_clk(i_clk));
Sub0000000002  u_000000057B_Sub0000000002(.i_data_1(A[175][1]), .i_data_2(B[175][1]), .o_data(mult_result_r[175][1]), .i_clk(i_clk));
Sub0000000002  u_000000057C_Sub0000000002(.i_data_1(B[175][1]), .i_data_2(C[175][1]), .o_data(mult_result_i[175][1]), .i_clk(i_clk));
Sub0000000002  u_000000057D_Sub0000000002(.i_data_1(A[175][2]), .i_data_2(B[175][2]), .o_data(mult_result_r[175][2]), .i_clk(i_clk));
Sub0000000002  u_000000057E_Sub0000000002(.i_data_1(B[175][2]), .i_data_2(C[175][2]), .o_data(mult_result_i[175][2]), .i_clk(i_clk));
Sub0000000002  u_000000057F_Sub0000000002(.i_data_1(A[175][3]), .i_data_2(B[175][3]), .o_data(mult_result_r[175][3]), .i_clk(i_clk));
Sub0000000002  u_0000000580_Sub0000000002(.i_data_1(B[175][3]), .i_data_2(C[175][3]), .o_data(mult_result_i[175][3]), .i_clk(i_clk));
Sub0000000002  u_0000000581_Sub0000000002(.i_data_1(A[176][0]), .i_data_2(B[176][0]), .o_data(mult_result_r[176][0]), .i_clk(i_clk));
Sub0000000002  u_0000000582_Sub0000000002(.i_data_1(B[176][0]), .i_data_2(C[176][0]), .o_data(mult_result_i[176][0]), .i_clk(i_clk));
Sub0000000002  u_0000000583_Sub0000000002(.i_data_1(A[176][1]), .i_data_2(B[176][1]), .o_data(mult_result_r[176][1]), .i_clk(i_clk));
Sub0000000002  u_0000000584_Sub0000000002(.i_data_1(B[176][1]), .i_data_2(C[176][1]), .o_data(mult_result_i[176][1]), .i_clk(i_clk));
Sub0000000002  u_0000000585_Sub0000000002(.i_data_1(A[176][2]), .i_data_2(B[176][2]), .o_data(mult_result_r[176][2]), .i_clk(i_clk));
Sub0000000002  u_0000000586_Sub0000000002(.i_data_1(B[176][2]), .i_data_2(C[176][2]), .o_data(mult_result_i[176][2]), .i_clk(i_clk));
Sub0000000002  u_0000000587_Sub0000000002(.i_data_1(A[176][3]), .i_data_2(B[176][3]), .o_data(mult_result_r[176][3]), .i_clk(i_clk));
Sub0000000002  u_0000000588_Sub0000000002(.i_data_1(B[176][3]), .i_data_2(C[176][3]), .o_data(mult_result_i[176][3]), .i_clk(i_clk));
Sub0000000002  u_0000000589_Sub0000000002(.i_data_1(A[177][0]), .i_data_2(B[177][0]), .o_data(mult_result_r[177][0]), .i_clk(i_clk));
Sub0000000002  u_000000058A_Sub0000000002(.i_data_1(B[177][0]), .i_data_2(C[177][0]), .o_data(mult_result_i[177][0]), .i_clk(i_clk));
Sub0000000002  u_000000058B_Sub0000000002(.i_data_1(A[177][1]), .i_data_2(B[177][1]), .o_data(mult_result_r[177][1]), .i_clk(i_clk));
Sub0000000002  u_000000058C_Sub0000000002(.i_data_1(B[177][1]), .i_data_2(C[177][1]), .o_data(mult_result_i[177][1]), .i_clk(i_clk));
Sub0000000002  u_000000058D_Sub0000000002(.i_data_1(A[177][2]), .i_data_2(B[177][2]), .o_data(mult_result_r[177][2]), .i_clk(i_clk));
Sub0000000002  u_000000058E_Sub0000000002(.i_data_1(B[177][2]), .i_data_2(C[177][2]), .o_data(mult_result_i[177][2]), .i_clk(i_clk));
Sub0000000002  u_000000058F_Sub0000000002(.i_data_1(A[177][3]), .i_data_2(B[177][3]), .o_data(mult_result_r[177][3]), .i_clk(i_clk));
Sub0000000002  u_0000000590_Sub0000000002(.i_data_1(B[177][3]), .i_data_2(C[177][3]), .o_data(mult_result_i[177][3]), .i_clk(i_clk));
Sub0000000002  u_0000000591_Sub0000000002(.i_data_1(A[178][0]), .i_data_2(B[178][0]), .o_data(mult_result_r[178][0]), .i_clk(i_clk));
Sub0000000002  u_0000000592_Sub0000000002(.i_data_1(B[178][0]), .i_data_2(C[178][0]), .o_data(mult_result_i[178][0]), .i_clk(i_clk));
Sub0000000002  u_0000000593_Sub0000000002(.i_data_1(A[178][1]), .i_data_2(B[178][1]), .o_data(mult_result_r[178][1]), .i_clk(i_clk));
Sub0000000002  u_0000000594_Sub0000000002(.i_data_1(B[178][1]), .i_data_2(C[178][1]), .o_data(mult_result_i[178][1]), .i_clk(i_clk));
Sub0000000002  u_0000000595_Sub0000000002(.i_data_1(A[178][2]), .i_data_2(B[178][2]), .o_data(mult_result_r[178][2]), .i_clk(i_clk));
Sub0000000002  u_0000000596_Sub0000000002(.i_data_1(B[178][2]), .i_data_2(C[178][2]), .o_data(mult_result_i[178][2]), .i_clk(i_clk));
Sub0000000002  u_0000000597_Sub0000000002(.i_data_1(A[178][3]), .i_data_2(B[178][3]), .o_data(mult_result_r[178][3]), .i_clk(i_clk));
Sub0000000002  u_0000000598_Sub0000000002(.i_data_1(B[178][3]), .i_data_2(C[178][3]), .o_data(mult_result_i[178][3]), .i_clk(i_clk));
Sub0000000002  u_0000000599_Sub0000000002(.i_data_1(A[179][0]), .i_data_2(B[179][0]), .o_data(mult_result_r[179][0]), .i_clk(i_clk));
Sub0000000002  u_000000059A_Sub0000000002(.i_data_1(B[179][0]), .i_data_2(C[179][0]), .o_data(mult_result_i[179][0]), .i_clk(i_clk));
Sub0000000002  u_000000059B_Sub0000000002(.i_data_1(A[179][1]), .i_data_2(B[179][1]), .o_data(mult_result_r[179][1]), .i_clk(i_clk));
Sub0000000002  u_000000059C_Sub0000000002(.i_data_1(B[179][1]), .i_data_2(C[179][1]), .o_data(mult_result_i[179][1]), .i_clk(i_clk));
Sub0000000002  u_000000059D_Sub0000000002(.i_data_1(A[179][2]), .i_data_2(B[179][2]), .o_data(mult_result_r[179][2]), .i_clk(i_clk));
Sub0000000002  u_000000059E_Sub0000000002(.i_data_1(B[179][2]), .i_data_2(C[179][2]), .o_data(mult_result_i[179][2]), .i_clk(i_clk));
Sub0000000002  u_000000059F_Sub0000000002(.i_data_1(A[179][3]), .i_data_2(B[179][3]), .o_data(mult_result_r[179][3]), .i_clk(i_clk));
Sub0000000002  u_00000005A0_Sub0000000002(.i_data_1(B[179][3]), .i_data_2(C[179][3]), .o_data(mult_result_i[179][3]), .i_clk(i_clk));
Sub0000000002  u_00000005A1_Sub0000000002(.i_data_1(A[180][0]), .i_data_2(B[180][0]), .o_data(mult_result_r[180][0]), .i_clk(i_clk));
Sub0000000002  u_00000005A2_Sub0000000002(.i_data_1(B[180][0]), .i_data_2(C[180][0]), .o_data(mult_result_i[180][0]), .i_clk(i_clk));
Sub0000000002  u_00000005A3_Sub0000000002(.i_data_1(A[180][1]), .i_data_2(B[180][1]), .o_data(mult_result_r[180][1]), .i_clk(i_clk));
Sub0000000002  u_00000005A4_Sub0000000002(.i_data_1(B[180][1]), .i_data_2(C[180][1]), .o_data(mult_result_i[180][1]), .i_clk(i_clk));
Sub0000000002  u_00000005A5_Sub0000000002(.i_data_1(A[180][2]), .i_data_2(B[180][2]), .o_data(mult_result_r[180][2]), .i_clk(i_clk));
Sub0000000002  u_00000005A6_Sub0000000002(.i_data_1(B[180][2]), .i_data_2(C[180][2]), .o_data(mult_result_i[180][2]), .i_clk(i_clk));
Sub0000000002  u_00000005A7_Sub0000000002(.i_data_1(A[180][3]), .i_data_2(B[180][3]), .o_data(mult_result_r[180][3]), .i_clk(i_clk));
Sub0000000002  u_00000005A8_Sub0000000002(.i_data_1(B[180][3]), .i_data_2(C[180][3]), .o_data(mult_result_i[180][3]), .i_clk(i_clk));
Sub0000000002  u_00000005A9_Sub0000000002(.i_data_1(A[181][0]), .i_data_2(B[181][0]), .o_data(mult_result_r[181][0]), .i_clk(i_clk));
Sub0000000002  u_00000005AA_Sub0000000002(.i_data_1(B[181][0]), .i_data_2(C[181][0]), .o_data(mult_result_i[181][0]), .i_clk(i_clk));
Sub0000000002  u_00000005AB_Sub0000000002(.i_data_1(A[181][1]), .i_data_2(B[181][1]), .o_data(mult_result_r[181][1]), .i_clk(i_clk));
Sub0000000002  u_00000005AC_Sub0000000002(.i_data_1(B[181][1]), .i_data_2(C[181][1]), .o_data(mult_result_i[181][1]), .i_clk(i_clk));
Sub0000000002  u_00000005AD_Sub0000000002(.i_data_1(A[181][2]), .i_data_2(B[181][2]), .o_data(mult_result_r[181][2]), .i_clk(i_clk));
Sub0000000002  u_00000005AE_Sub0000000002(.i_data_1(B[181][2]), .i_data_2(C[181][2]), .o_data(mult_result_i[181][2]), .i_clk(i_clk));
Sub0000000002  u_00000005AF_Sub0000000002(.i_data_1(A[181][3]), .i_data_2(B[181][3]), .o_data(mult_result_r[181][3]), .i_clk(i_clk));
Sub0000000002  u_00000005B0_Sub0000000002(.i_data_1(B[181][3]), .i_data_2(C[181][3]), .o_data(mult_result_i[181][3]), .i_clk(i_clk));
Sub0000000002  u_00000005B1_Sub0000000002(.i_data_1(A[182][0]), .i_data_2(B[182][0]), .o_data(mult_result_r[182][0]), .i_clk(i_clk));
Sub0000000002  u_00000005B2_Sub0000000002(.i_data_1(B[182][0]), .i_data_2(C[182][0]), .o_data(mult_result_i[182][0]), .i_clk(i_clk));
Sub0000000002  u_00000005B3_Sub0000000002(.i_data_1(A[182][1]), .i_data_2(B[182][1]), .o_data(mult_result_r[182][1]), .i_clk(i_clk));
Sub0000000002  u_00000005B4_Sub0000000002(.i_data_1(B[182][1]), .i_data_2(C[182][1]), .o_data(mult_result_i[182][1]), .i_clk(i_clk));
Sub0000000002  u_00000005B5_Sub0000000002(.i_data_1(A[182][2]), .i_data_2(B[182][2]), .o_data(mult_result_r[182][2]), .i_clk(i_clk));
Sub0000000002  u_00000005B6_Sub0000000002(.i_data_1(B[182][2]), .i_data_2(C[182][2]), .o_data(mult_result_i[182][2]), .i_clk(i_clk));
Sub0000000002  u_00000005B7_Sub0000000002(.i_data_1(A[182][3]), .i_data_2(B[182][3]), .o_data(mult_result_r[182][3]), .i_clk(i_clk));
Sub0000000002  u_00000005B8_Sub0000000002(.i_data_1(B[182][3]), .i_data_2(C[182][3]), .o_data(mult_result_i[182][3]), .i_clk(i_clk));
Sub0000000002  u_00000005B9_Sub0000000002(.i_data_1(A[183][0]), .i_data_2(B[183][0]), .o_data(mult_result_r[183][0]), .i_clk(i_clk));
Sub0000000002  u_00000005BA_Sub0000000002(.i_data_1(B[183][0]), .i_data_2(C[183][0]), .o_data(mult_result_i[183][0]), .i_clk(i_clk));
Sub0000000002  u_00000005BB_Sub0000000002(.i_data_1(A[183][1]), .i_data_2(B[183][1]), .o_data(mult_result_r[183][1]), .i_clk(i_clk));
Sub0000000002  u_00000005BC_Sub0000000002(.i_data_1(B[183][1]), .i_data_2(C[183][1]), .o_data(mult_result_i[183][1]), .i_clk(i_clk));
Sub0000000002  u_00000005BD_Sub0000000002(.i_data_1(A[183][2]), .i_data_2(B[183][2]), .o_data(mult_result_r[183][2]), .i_clk(i_clk));
Sub0000000002  u_00000005BE_Sub0000000002(.i_data_1(B[183][2]), .i_data_2(C[183][2]), .o_data(mult_result_i[183][2]), .i_clk(i_clk));
Sub0000000002  u_00000005BF_Sub0000000002(.i_data_1(A[183][3]), .i_data_2(B[183][3]), .o_data(mult_result_r[183][3]), .i_clk(i_clk));
Sub0000000002  u_00000005C0_Sub0000000002(.i_data_1(B[183][3]), .i_data_2(C[183][3]), .o_data(mult_result_i[183][3]), .i_clk(i_clk));
Sub0000000002  u_00000005C1_Sub0000000002(.i_data_1(A[184][0]), .i_data_2(B[184][0]), .o_data(mult_result_r[184][0]), .i_clk(i_clk));
Sub0000000002  u_00000005C2_Sub0000000002(.i_data_1(B[184][0]), .i_data_2(C[184][0]), .o_data(mult_result_i[184][0]), .i_clk(i_clk));
Sub0000000002  u_00000005C3_Sub0000000002(.i_data_1(A[184][1]), .i_data_2(B[184][1]), .o_data(mult_result_r[184][1]), .i_clk(i_clk));
Sub0000000002  u_00000005C4_Sub0000000002(.i_data_1(B[184][1]), .i_data_2(C[184][1]), .o_data(mult_result_i[184][1]), .i_clk(i_clk));
Sub0000000002  u_00000005C5_Sub0000000002(.i_data_1(A[184][2]), .i_data_2(B[184][2]), .o_data(mult_result_r[184][2]), .i_clk(i_clk));
Sub0000000002  u_00000005C6_Sub0000000002(.i_data_1(B[184][2]), .i_data_2(C[184][2]), .o_data(mult_result_i[184][2]), .i_clk(i_clk));
Sub0000000002  u_00000005C7_Sub0000000002(.i_data_1(A[184][3]), .i_data_2(B[184][3]), .o_data(mult_result_r[184][3]), .i_clk(i_clk));
Sub0000000002  u_00000005C8_Sub0000000002(.i_data_1(B[184][3]), .i_data_2(C[184][3]), .o_data(mult_result_i[184][3]), .i_clk(i_clk));
Sub0000000002  u_00000005C9_Sub0000000002(.i_data_1(A[185][0]), .i_data_2(B[185][0]), .o_data(mult_result_r[185][0]), .i_clk(i_clk));
Sub0000000002  u_00000005CA_Sub0000000002(.i_data_1(B[185][0]), .i_data_2(C[185][0]), .o_data(mult_result_i[185][0]), .i_clk(i_clk));
Sub0000000002  u_00000005CB_Sub0000000002(.i_data_1(A[185][1]), .i_data_2(B[185][1]), .o_data(mult_result_r[185][1]), .i_clk(i_clk));
Sub0000000002  u_00000005CC_Sub0000000002(.i_data_1(B[185][1]), .i_data_2(C[185][1]), .o_data(mult_result_i[185][1]), .i_clk(i_clk));
Sub0000000002  u_00000005CD_Sub0000000002(.i_data_1(A[185][2]), .i_data_2(B[185][2]), .o_data(mult_result_r[185][2]), .i_clk(i_clk));
Sub0000000002  u_00000005CE_Sub0000000002(.i_data_1(B[185][2]), .i_data_2(C[185][2]), .o_data(mult_result_i[185][2]), .i_clk(i_clk));
Sub0000000002  u_00000005CF_Sub0000000002(.i_data_1(A[185][3]), .i_data_2(B[185][3]), .o_data(mult_result_r[185][3]), .i_clk(i_clk));
Sub0000000002  u_00000005D0_Sub0000000002(.i_data_1(B[185][3]), .i_data_2(C[185][3]), .o_data(mult_result_i[185][3]), .i_clk(i_clk));
Sub0000000002  u_00000005D1_Sub0000000002(.i_data_1(A[186][0]), .i_data_2(B[186][0]), .o_data(mult_result_r[186][0]), .i_clk(i_clk));
Sub0000000002  u_00000005D2_Sub0000000002(.i_data_1(B[186][0]), .i_data_2(C[186][0]), .o_data(mult_result_i[186][0]), .i_clk(i_clk));
Sub0000000002  u_00000005D3_Sub0000000002(.i_data_1(A[186][1]), .i_data_2(B[186][1]), .o_data(mult_result_r[186][1]), .i_clk(i_clk));
Sub0000000002  u_00000005D4_Sub0000000002(.i_data_1(B[186][1]), .i_data_2(C[186][1]), .o_data(mult_result_i[186][1]), .i_clk(i_clk));
Sub0000000002  u_00000005D5_Sub0000000002(.i_data_1(A[186][2]), .i_data_2(B[186][2]), .o_data(mult_result_r[186][2]), .i_clk(i_clk));
Sub0000000002  u_00000005D6_Sub0000000002(.i_data_1(B[186][2]), .i_data_2(C[186][2]), .o_data(mult_result_i[186][2]), .i_clk(i_clk));
Sub0000000002  u_00000005D7_Sub0000000002(.i_data_1(A[186][3]), .i_data_2(B[186][3]), .o_data(mult_result_r[186][3]), .i_clk(i_clk));
Sub0000000002  u_00000005D8_Sub0000000002(.i_data_1(B[186][3]), .i_data_2(C[186][3]), .o_data(mult_result_i[186][3]), .i_clk(i_clk));
Sub0000000002  u_00000005D9_Sub0000000002(.i_data_1(A[187][0]), .i_data_2(B[187][0]), .o_data(mult_result_r[187][0]), .i_clk(i_clk));
Sub0000000002  u_00000005DA_Sub0000000002(.i_data_1(B[187][0]), .i_data_2(C[187][0]), .o_data(mult_result_i[187][0]), .i_clk(i_clk));
Sub0000000002  u_00000005DB_Sub0000000002(.i_data_1(A[187][1]), .i_data_2(B[187][1]), .o_data(mult_result_r[187][1]), .i_clk(i_clk));
Sub0000000002  u_00000005DC_Sub0000000002(.i_data_1(B[187][1]), .i_data_2(C[187][1]), .o_data(mult_result_i[187][1]), .i_clk(i_clk));
Sub0000000002  u_00000005DD_Sub0000000002(.i_data_1(A[187][2]), .i_data_2(B[187][2]), .o_data(mult_result_r[187][2]), .i_clk(i_clk));
Sub0000000002  u_00000005DE_Sub0000000002(.i_data_1(B[187][2]), .i_data_2(C[187][2]), .o_data(mult_result_i[187][2]), .i_clk(i_clk));
Sub0000000002  u_00000005DF_Sub0000000002(.i_data_1(A[187][3]), .i_data_2(B[187][3]), .o_data(mult_result_r[187][3]), .i_clk(i_clk));
Sub0000000002  u_00000005E0_Sub0000000002(.i_data_1(B[187][3]), .i_data_2(C[187][3]), .o_data(mult_result_i[187][3]), .i_clk(i_clk));
Sub0000000002  u_00000005E1_Sub0000000002(.i_data_1(A[188][0]), .i_data_2(B[188][0]), .o_data(mult_result_r[188][0]), .i_clk(i_clk));
Sub0000000002  u_00000005E2_Sub0000000002(.i_data_1(B[188][0]), .i_data_2(C[188][0]), .o_data(mult_result_i[188][0]), .i_clk(i_clk));
Sub0000000002  u_00000005E3_Sub0000000002(.i_data_1(A[188][1]), .i_data_2(B[188][1]), .o_data(mult_result_r[188][1]), .i_clk(i_clk));
Sub0000000002  u_00000005E4_Sub0000000002(.i_data_1(B[188][1]), .i_data_2(C[188][1]), .o_data(mult_result_i[188][1]), .i_clk(i_clk));
Sub0000000002  u_00000005E5_Sub0000000002(.i_data_1(A[188][2]), .i_data_2(B[188][2]), .o_data(mult_result_r[188][2]), .i_clk(i_clk));
Sub0000000002  u_00000005E6_Sub0000000002(.i_data_1(B[188][2]), .i_data_2(C[188][2]), .o_data(mult_result_i[188][2]), .i_clk(i_clk));
Sub0000000002  u_00000005E7_Sub0000000002(.i_data_1(A[188][3]), .i_data_2(B[188][3]), .o_data(mult_result_r[188][3]), .i_clk(i_clk));
Sub0000000002  u_00000005E8_Sub0000000002(.i_data_1(B[188][3]), .i_data_2(C[188][3]), .o_data(mult_result_i[188][3]), .i_clk(i_clk));
Sub0000000002  u_00000005E9_Sub0000000002(.i_data_1(A[189][0]), .i_data_2(B[189][0]), .o_data(mult_result_r[189][0]), .i_clk(i_clk));
Sub0000000002  u_00000005EA_Sub0000000002(.i_data_1(B[189][0]), .i_data_2(C[189][0]), .o_data(mult_result_i[189][0]), .i_clk(i_clk));
Sub0000000002  u_00000005EB_Sub0000000002(.i_data_1(A[189][1]), .i_data_2(B[189][1]), .o_data(mult_result_r[189][1]), .i_clk(i_clk));
Sub0000000002  u_00000005EC_Sub0000000002(.i_data_1(B[189][1]), .i_data_2(C[189][1]), .o_data(mult_result_i[189][1]), .i_clk(i_clk));
Sub0000000002  u_00000005ED_Sub0000000002(.i_data_1(A[189][2]), .i_data_2(B[189][2]), .o_data(mult_result_r[189][2]), .i_clk(i_clk));
Sub0000000002  u_00000005EE_Sub0000000002(.i_data_1(B[189][2]), .i_data_2(C[189][2]), .o_data(mult_result_i[189][2]), .i_clk(i_clk));
Sub0000000002  u_00000005EF_Sub0000000002(.i_data_1(A[189][3]), .i_data_2(B[189][3]), .o_data(mult_result_r[189][3]), .i_clk(i_clk));
Sub0000000002  u_00000005F0_Sub0000000002(.i_data_1(B[189][3]), .i_data_2(C[189][3]), .o_data(mult_result_i[189][3]), .i_clk(i_clk));
Sub0000000002  u_00000005F1_Sub0000000002(.i_data_1(A[190][0]), .i_data_2(B[190][0]), .o_data(mult_result_r[190][0]), .i_clk(i_clk));
Sub0000000002  u_00000005F2_Sub0000000002(.i_data_1(B[190][0]), .i_data_2(C[190][0]), .o_data(mult_result_i[190][0]), .i_clk(i_clk));
Sub0000000002  u_00000005F3_Sub0000000002(.i_data_1(A[190][1]), .i_data_2(B[190][1]), .o_data(mult_result_r[190][1]), .i_clk(i_clk));
Sub0000000002  u_00000005F4_Sub0000000002(.i_data_1(B[190][1]), .i_data_2(C[190][1]), .o_data(mult_result_i[190][1]), .i_clk(i_clk));
Sub0000000002  u_00000005F5_Sub0000000002(.i_data_1(A[190][2]), .i_data_2(B[190][2]), .o_data(mult_result_r[190][2]), .i_clk(i_clk));
Sub0000000002  u_00000005F6_Sub0000000002(.i_data_1(B[190][2]), .i_data_2(C[190][2]), .o_data(mult_result_i[190][2]), .i_clk(i_clk));
Sub0000000002  u_00000005F7_Sub0000000002(.i_data_1(A[190][3]), .i_data_2(B[190][3]), .o_data(mult_result_r[190][3]), .i_clk(i_clk));
Sub0000000002  u_00000005F8_Sub0000000002(.i_data_1(B[190][3]), .i_data_2(C[190][3]), .o_data(mult_result_i[190][3]), .i_clk(i_clk));
Sub0000000002  u_00000005F9_Sub0000000002(.i_data_1(A[191][0]), .i_data_2(B[191][0]), .o_data(mult_result_r[191][0]), .i_clk(i_clk));
Sub0000000002  u_00000005FA_Sub0000000002(.i_data_1(B[191][0]), .i_data_2(C[191][0]), .o_data(mult_result_i[191][0]), .i_clk(i_clk));
Sub0000000002  u_00000005FB_Sub0000000002(.i_data_1(A[191][1]), .i_data_2(B[191][1]), .o_data(mult_result_r[191][1]), .i_clk(i_clk));
Sub0000000002  u_00000005FC_Sub0000000002(.i_data_1(B[191][1]), .i_data_2(C[191][1]), .o_data(mult_result_i[191][1]), .i_clk(i_clk));
Sub0000000002  u_00000005FD_Sub0000000002(.i_data_1(A[191][2]), .i_data_2(B[191][2]), .o_data(mult_result_r[191][2]), .i_clk(i_clk));
Sub0000000002  u_00000005FE_Sub0000000002(.i_data_1(B[191][2]), .i_data_2(C[191][2]), .o_data(mult_result_i[191][2]), .i_clk(i_clk));
Sub0000000002  u_00000005FF_Sub0000000002(.i_data_1(A[191][3]), .i_data_2(B[191][3]), .o_data(mult_result_r[191][3]), .i_clk(i_clk));
Sub0000000002  u_0000000600_Sub0000000002(.i_data_1(B[191][3]), .i_data_2(C[191][3]), .o_data(mult_result_i[191][3]), .i_clk(i_clk));
Sub0000000002  u_0000000601_Sub0000000002(.i_data_1(A[192][0]), .i_data_2(B[192][0]), .o_data(mult_result_r[192][0]), .i_clk(i_clk));
Sub0000000002  u_0000000602_Sub0000000002(.i_data_1(B[192][0]), .i_data_2(C[192][0]), .o_data(mult_result_i[192][0]), .i_clk(i_clk));
Sub0000000002  u_0000000603_Sub0000000002(.i_data_1(A[192][1]), .i_data_2(B[192][1]), .o_data(mult_result_r[192][1]), .i_clk(i_clk));
Sub0000000002  u_0000000604_Sub0000000002(.i_data_1(B[192][1]), .i_data_2(C[192][1]), .o_data(mult_result_i[192][1]), .i_clk(i_clk));
Sub0000000002  u_0000000605_Sub0000000002(.i_data_1(A[192][2]), .i_data_2(B[192][2]), .o_data(mult_result_r[192][2]), .i_clk(i_clk));
Sub0000000002  u_0000000606_Sub0000000002(.i_data_1(B[192][2]), .i_data_2(C[192][2]), .o_data(mult_result_i[192][2]), .i_clk(i_clk));
Sub0000000002  u_0000000607_Sub0000000002(.i_data_1(A[192][3]), .i_data_2(B[192][3]), .o_data(mult_result_r[192][3]), .i_clk(i_clk));
Sub0000000002  u_0000000608_Sub0000000002(.i_data_1(B[192][3]), .i_data_2(C[192][3]), .o_data(mult_result_i[192][3]), .i_clk(i_clk));
Sub0000000002  u_0000000609_Sub0000000002(.i_data_1(A[193][0]), .i_data_2(B[193][0]), .o_data(mult_result_r[193][0]), .i_clk(i_clk));
Sub0000000002  u_000000060A_Sub0000000002(.i_data_1(B[193][0]), .i_data_2(C[193][0]), .o_data(mult_result_i[193][0]), .i_clk(i_clk));
Sub0000000002  u_000000060B_Sub0000000002(.i_data_1(A[193][1]), .i_data_2(B[193][1]), .o_data(mult_result_r[193][1]), .i_clk(i_clk));
Sub0000000002  u_000000060C_Sub0000000002(.i_data_1(B[193][1]), .i_data_2(C[193][1]), .o_data(mult_result_i[193][1]), .i_clk(i_clk));
Sub0000000002  u_000000060D_Sub0000000002(.i_data_1(A[193][2]), .i_data_2(B[193][2]), .o_data(mult_result_r[193][2]), .i_clk(i_clk));
Sub0000000002  u_000000060E_Sub0000000002(.i_data_1(B[193][2]), .i_data_2(C[193][2]), .o_data(mult_result_i[193][2]), .i_clk(i_clk));
Sub0000000002  u_000000060F_Sub0000000002(.i_data_1(A[193][3]), .i_data_2(B[193][3]), .o_data(mult_result_r[193][3]), .i_clk(i_clk));
Sub0000000002  u_0000000610_Sub0000000002(.i_data_1(B[193][3]), .i_data_2(C[193][3]), .o_data(mult_result_i[193][3]), .i_clk(i_clk));
Sub0000000002  u_0000000611_Sub0000000002(.i_data_1(A[194][0]), .i_data_2(B[194][0]), .o_data(mult_result_r[194][0]), .i_clk(i_clk));
Sub0000000002  u_0000000612_Sub0000000002(.i_data_1(B[194][0]), .i_data_2(C[194][0]), .o_data(mult_result_i[194][0]), .i_clk(i_clk));
Sub0000000002  u_0000000613_Sub0000000002(.i_data_1(A[194][1]), .i_data_2(B[194][1]), .o_data(mult_result_r[194][1]), .i_clk(i_clk));
Sub0000000002  u_0000000614_Sub0000000002(.i_data_1(B[194][1]), .i_data_2(C[194][1]), .o_data(mult_result_i[194][1]), .i_clk(i_clk));
Sub0000000002  u_0000000615_Sub0000000002(.i_data_1(A[194][2]), .i_data_2(B[194][2]), .o_data(mult_result_r[194][2]), .i_clk(i_clk));
Sub0000000002  u_0000000616_Sub0000000002(.i_data_1(B[194][2]), .i_data_2(C[194][2]), .o_data(mult_result_i[194][2]), .i_clk(i_clk));
Sub0000000002  u_0000000617_Sub0000000002(.i_data_1(A[194][3]), .i_data_2(B[194][3]), .o_data(mult_result_r[194][3]), .i_clk(i_clk));
Sub0000000002  u_0000000618_Sub0000000002(.i_data_1(B[194][3]), .i_data_2(C[194][3]), .o_data(mult_result_i[194][3]), .i_clk(i_clk));
Sub0000000002  u_0000000619_Sub0000000002(.i_data_1(A[195][0]), .i_data_2(B[195][0]), .o_data(mult_result_r[195][0]), .i_clk(i_clk));
Sub0000000002  u_000000061A_Sub0000000002(.i_data_1(B[195][0]), .i_data_2(C[195][0]), .o_data(mult_result_i[195][0]), .i_clk(i_clk));
Sub0000000002  u_000000061B_Sub0000000002(.i_data_1(A[195][1]), .i_data_2(B[195][1]), .o_data(mult_result_r[195][1]), .i_clk(i_clk));
Sub0000000002  u_000000061C_Sub0000000002(.i_data_1(B[195][1]), .i_data_2(C[195][1]), .o_data(mult_result_i[195][1]), .i_clk(i_clk));
Sub0000000002  u_000000061D_Sub0000000002(.i_data_1(A[195][2]), .i_data_2(B[195][2]), .o_data(mult_result_r[195][2]), .i_clk(i_clk));
Sub0000000002  u_000000061E_Sub0000000002(.i_data_1(B[195][2]), .i_data_2(C[195][2]), .o_data(mult_result_i[195][2]), .i_clk(i_clk));
Sub0000000002  u_000000061F_Sub0000000002(.i_data_1(A[195][3]), .i_data_2(B[195][3]), .o_data(mult_result_r[195][3]), .i_clk(i_clk));
Sub0000000002  u_0000000620_Sub0000000002(.i_data_1(B[195][3]), .i_data_2(C[195][3]), .o_data(mult_result_i[195][3]), .i_clk(i_clk));
Sub0000000002  u_0000000621_Sub0000000002(.i_data_1(A[196][0]), .i_data_2(B[196][0]), .o_data(mult_result_r[196][0]), .i_clk(i_clk));
Sub0000000002  u_0000000622_Sub0000000002(.i_data_1(B[196][0]), .i_data_2(C[196][0]), .o_data(mult_result_i[196][0]), .i_clk(i_clk));
Sub0000000002  u_0000000623_Sub0000000002(.i_data_1(A[196][1]), .i_data_2(B[196][1]), .o_data(mult_result_r[196][1]), .i_clk(i_clk));
Sub0000000002  u_0000000624_Sub0000000002(.i_data_1(B[196][1]), .i_data_2(C[196][1]), .o_data(mult_result_i[196][1]), .i_clk(i_clk));
Sub0000000002  u_0000000625_Sub0000000002(.i_data_1(A[196][2]), .i_data_2(B[196][2]), .o_data(mult_result_r[196][2]), .i_clk(i_clk));
Sub0000000002  u_0000000626_Sub0000000002(.i_data_1(B[196][2]), .i_data_2(C[196][2]), .o_data(mult_result_i[196][2]), .i_clk(i_clk));
Sub0000000002  u_0000000627_Sub0000000002(.i_data_1(A[196][3]), .i_data_2(B[196][3]), .o_data(mult_result_r[196][3]), .i_clk(i_clk));
Sub0000000002  u_0000000628_Sub0000000002(.i_data_1(B[196][3]), .i_data_2(C[196][3]), .o_data(mult_result_i[196][3]), .i_clk(i_clk));
Sub0000000002  u_0000000629_Sub0000000002(.i_data_1(A[197][0]), .i_data_2(B[197][0]), .o_data(mult_result_r[197][0]), .i_clk(i_clk));
Sub0000000002  u_000000062A_Sub0000000002(.i_data_1(B[197][0]), .i_data_2(C[197][0]), .o_data(mult_result_i[197][0]), .i_clk(i_clk));
Sub0000000002  u_000000062B_Sub0000000002(.i_data_1(A[197][1]), .i_data_2(B[197][1]), .o_data(mult_result_r[197][1]), .i_clk(i_clk));
Sub0000000002  u_000000062C_Sub0000000002(.i_data_1(B[197][1]), .i_data_2(C[197][1]), .o_data(mult_result_i[197][1]), .i_clk(i_clk));
Sub0000000002  u_000000062D_Sub0000000002(.i_data_1(A[197][2]), .i_data_2(B[197][2]), .o_data(mult_result_r[197][2]), .i_clk(i_clk));
Sub0000000002  u_000000062E_Sub0000000002(.i_data_1(B[197][2]), .i_data_2(C[197][2]), .o_data(mult_result_i[197][2]), .i_clk(i_clk));
Sub0000000002  u_000000062F_Sub0000000002(.i_data_1(A[197][3]), .i_data_2(B[197][3]), .o_data(mult_result_r[197][3]), .i_clk(i_clk));
Sub0000000002  u_0000000630_Sub0000000002(.i_data_1(B[197][3]), .i_data_2(C[197][3]), .o_data(mult_result_i[197][3]), .i_clk(i_clk));
Sub0000000002  u_0000000631_Sub0000000002(.i_data_1(A[198][0]), .i_data_2(B[198][0]), .o_data(mult_result_r[198][0]), .i_clk(i_clk));
Sub0000000002  u_0000000632_Sub0000000002(.i_data_1(B[198][0]), .i_data_2(C[198][0]), .o_data(mult_result_i[198][0]), .i_clk(i_clk));
Sub0000000002  u_0000000633_Sub0000000002(.i_data_1(A[198][1]), .i_data_2(B[198][1]), .o_data(mult_result_r[198][1]), .i_clk(i_clk));
Sub0000000002  u_0000000634_Sub0000000002(.i_data_1(B[198][1]), .i_data_2(C[198][1]), .o_data(mult_result_i[198][1]), .i_clk(i_clk));
Sub0000000002  u_0000000635_Sub0000000002(.i_data_1(A[198][2]), .i_data_2(B[198][2]), .o_data(mult_result_r[198][2]), .i_clk(i_clk));
Sub0000000002  u_0000000636_Sub0000000002(.i_data_1(B[198][2]), .i_data_2(C[198][2]), .o_data(mult_result_i[198][2]), .i_clk(i_clk));
Sub0000000002  u_0000000637_Sub0000000002(.i_data_1(A[198][3]), .i_data_2(B[198][3]), .o_data(mult_result_r[198][3]), .i_clk(i_clk));
Sub0000000002  u_0000000638_Sub0000000002(.i_data_1(B[198][3]), .i_data_2(C[198][3]), .o_data(mult_result_i[198][3]), .i_clk(i_clk));
Sub0000000002  u_0000000639_Sub0000000002(.i_data_1(A[199][0]), .i_data_2(B[199][0]), .o_data(mult_result_r[199][0]), .i_clk(i_clk));
Sub0000000002  u_000000063A_Sub0000000002(.i_data_1(B[199][0]), .i_data_2(C[199][0]), .o_data(mult_result_i[199][0]), .i_clk(i_clk));
Sub0000000002  u_000000063B_Sub0000000002(.i_data_1(A[199][1]), .i_data_2(B[199][1]), .o_data(mult_result_r[199][1]), .i_clk(i_clk));
Sub0000000002  u_000000063C_Sub0000000002(.i_data_1(B[199][1]), .i_data_2(C[199][1]), .o_data(mult_result_i[199][1]), .i_clk(i_clk));
Sub0000000002  u_000000063D_Sub0000000002(.i_data_1(A[199][2]), .i_data_2(B[199][2]), .o_data(mult_result_r[199][2]), .i_clk(i_clk));
Sub0000000002  u_000000063E_Sub0000000002(.i_data_1(B[199][2]), .i_data_2(C[199][2]), .o_data(mult_result_i[199][2]), .i_clk(i_clk));
Sub0000000002  u_000000063F_Sub0000000002(.i_data_1(A[199][3]), .i_data_2(B[199][3]), .o_data(mult_result_r[199][3]), .i_clk(i_clk));
Sub0000000002  u_0000000640_Sub0000000002(.i_data_1(B[199][3]), .i_data_2(C[199][3]), .o_data(mult_result_i[199][3]), .i_clk(i_clk));
Sub0000000002  u_0000000641_Sub0000000002(.i_data_1(A[200][0]), .i_data_2(B[200][0]), .o_data(mult_result_r[200][0]), .i_clk(i_clk));
Sub0000000002  u_0000000642_Sub0000000002(.i_data_1(B[200][0]), .i_data_2(C[200][0]), .o_data(mult_result_i[200][0]), .i_clk(i_clk));
Sub0000000002  u_0000000643_Sub0000000002(.i_data_1(A[200][1]), .i_data_2(B[200][1]), .o_data(mult_result_r[200][1]), .i_clk(i_clk));
Sub0000000002  u_0000000644_Sub0000000002(.i_data_1(B[200][1]), .i_data_2(C[200][1]), .o_data(mult_result_i[200][1]), .i_clk(i_clk));
Sub0000000002  u_0000000645_Sub0000000002(.i_data_1(A[200][2]), .i_data_2(B[200][2]), .o_data(mult_result_r[200][2]), .i_clk(i_clk));
Sub0000000002  u_0000000646_Sub0000000002(.i_data_1(B[200][2]), .i_data_2(C[200][2]), .o_data(mult_result_i[200][2]), .i_clk(i_clk));
Sub0000000002  u_0000000647_Sub0000000002(.i_data_1(A[200][3]), .i_data_2(B[200][3]), .o_data(mult_result_r[200][3]), .i_clk(i_clk));
Sub0000000002  u_0000000648_Sub0000000002(.i_data_1(B[200][3]), .i_data_2(C[200][3]), .o_data(mult_result_i[200][3]), .i_clk(i_clk));
Sub0000000002  u_0000000649_Sub0000000002(.i_data_1(A[201][0]), .i_data_2(B[201][0]), .o_data(mult_result_r[201][0]), .i_clk(i_clk));
Sub0000000002  u_000000064A_Sub0000000002(.i_data_1(B[201][0]), .i_data_2(C[201][0]), .o_data(mult_result_i[201][0]), .i_clk(i_clk));
Sub0000000002  u_000000064B_Sub0000000002(.i_data_1(A[201][1]), .i_data_2(B[201][1]), .o_data(mult_result_r[201][1]), .i_clk(i_clk));
Sub0000000002  u_000000064C_Sub0000000002(.i_data_1(B[201][1]), .i_data_2(C[201][1]), .o_data(mult_result_i[201][1]), .i_clk(i_clk));
Sub0000000002  u_000000064D_Sub0000000002(.i_data_1(A[201][2]), .i_data_2(B[201][2]), .o_data(mult_result_r[201][2]), .i_clk(i_clk));
Sub0000000002  u_000000064E_Sub0000000002(.i_data_1(B[201][2]), .i_data_2(C[201][2]), .o_data(mult_result_i[201][2]), .i_clk(i_clk));
Sub0000000002  u_000000064F_Sub0000000002(.i_data_1(A[201][3]), .i_data_2(B[201][3]), .o_data(mult_result_r[201][3]), .i_clk(i_clk));
Sub0000000002  u_0000000650_Sub0000000002(.i_data_1(B[201][3]), .i_data_2(C[201][3]), .o_data(mult_result_i[201][3]), .i_clk(i_clk));
Sub0000000002  u_0000000651_Sub0000000002(.i_data_1(A[202][0]), .i_data_2(B[202][0]), .o_data(mult_result_r[202][0]), .i_clk(i_clk));
Sub0000000002  u_0000000652_Sub0000000002(.i_data_1(B[202][0]), .i_data_2(C[202][0]), .o_data(mult_result_i[202][0]), .i_clk(i_clk));
Sub0000000002  u_0000000653_Sub0000000002(.i_data_1(A[202][1]), .i_data_2(B[202][1]), .o_data(mult_result_r[202][1]), .i_clk(i_clk));
Sub0000000002  u_0000000654_Sub0000000002(.i_data_1(B[202][1]), .i_data_2(C[202][1]), .o_data(mult_result_i[202][1]), .i_clk(i_clk));
Sub0000000002  u_0000000655_Sub0000000002(.i_data_1(A[202][2]), .i_data_2(B[202][2]), .o_data(mult_result_r[202][2]), .i_clk(i_clk));
Sub0000000002  u_0000000656_Sub0000000002(.i_data_1(B[202][2]), .i_data_2(C[202][2]), .o_data(mult_result_i[202][2]), .i_clk(i_clk));
Sub0000000002  u_0000000657_Sub0000000002(.i_data_1(A[202][3]), .i_data_2(B[202][3]), .o_data(mult_result_r[202][3]), .i_clk(i_clk));
Sub0000000002  u_0000000658_Sub0000000002(.i_data_1(B[202][3]), .i_data_2(C[202][3]), .o_data(mult_result_i[202][3]), .i_clk(i_clk));
Sub0000000002  u_0000000659_Sub0000000002(.i_data_1(A[203][0]), .i_data_2(B[203][0]), .o_data(mult_result_r[203][0]), .i_clk(i_clk));
Sub0000000002  u_000000065A_Sub0000000002(.i_data_1(B[203][0]), .i_data_2(C[203][0]), .o_data(mult_result_i[203][0]), .i_clk(i_clk));
Sub0000000002  u_000000065B_Sub0000000002(.i_data_1(A[203][1]), .i_data_2(B[203][1]), .o_data(mult_result_r[203][1]), .i_clk(i_clk));
Sub0000000002  u_000000065C_Sub0000000002(.i_data_1(B[203][1]), .i_data_2(C[203][1]), .o_data(mult_result_i[203][1]), .i_clk(i_clk));
Sub0000000002  u_000000065D_Sub0000000002(.i_data_1(A[203][2]), .i_data_2(B[203][2]), .o_data(mult_result_r[203][2]), .i_clk(i_clk));
Sub0000000002  u_000000065E_Sub0000000002(.i_data_1(B[203][2]), .i_data_2(C[203][2]), .o_data(mult_result_i[203][2]), .i_clk(i_clk));
Sub0000000002  u_000000065F_Sub0000000002(.i_data_1(A[203][3]), .i_data_2(B[203][3]), .o_data(mult_result_r[203][3]), .i_clk(i_clk));
Sub0000000002  u_0000000660_Sub0000000002(.i_data_1(B[203][3]), .i_data_2(C[203][3]), .o_data(mult_result_i[203][3]), .i_clk(i_clk));
Sub0000000002  u_0000000661_Sub0000000002(.i_data_1(A[204][0]), .i_data_2(B[204][0]), .o_data(mult_result_r[204][0]), .i_clk(i_clk));
Sub0000000002  u_0000000662_Sub0000000002(.i_data_1(B[204][0]), .i_data_2(C[204][0]), .o_data(mult_result_i[204][0]), .i_clk(i_clk));
Sub0000000002  u_0000000663_Sub0000000002(.i_data_1(A[204][1]), .i_data_2(B[204][1]), .o_data(mult_result_r[204][1]), .i_clk(i_clk));
Sub0000000002  u_0000000664_Sub0000000002(.i_data_1(B[204][1]), .i_data_2(C[204][1]), .o_data(mult_result_i[204][1]), .i_clk(i_clk));
Sub0000000002  u_0000000665_Sub0000000002(.i_data_1(A[204][2]), .i_data_2(B[204][2]), .o_data(mult_result_r[204][2]), .i_clk(i_clk));
Sub0000000002  u_0000000666_Sub0000000002(.i_data_1(B[204][2]), .i_data_2(C[204][2]), .o_data(mult_result_i[204][2]), .i_clk(i_clk));
Sub0000000002  u_0000000667_Sub0000000002(.i_data_1(A[204][3]), .i_data_2(B[204][3]), .o_data(mult_result_r[204][3]), .i_clk(i_clk));
Sub0000000002  u_0000000668_Sub0000000002(.i_data_1(B[204][3]), .i_data_2(C[204][3]), .o_data(mult_result_i[204][3]), .i_clk(i_clk));
Sub0000000002  u_0000000669_Sub0000000002(.i_data_1(A[205][0]), .i_data_2(B[205][0]), .o_data(mult_result_r[205][0]), .i_clk(i_clk));
Sub0000000002  u_000000066A_Sub0000000002(.i_data_1(B[205][0]), .i_data_2(C[205][0]), .o_data(mult_result_i[205][0]), .i_clk(i_clk));
Sub0000000002  u_000000066B_Sub0000000002(.i_data_1(A[205][1]), .i_data_2(B[205][1]), .o_data(mult_result_r[205][1]), .i_clk(i_clk));
Sub0000000002  u_000000066C_Sub0000000002(.i_data_1(B[205][1]), .i_data_2(C[205][1]), .o_data(mult_result_i[205][1]), .i_clk(i_clk));
Sub0000000002  u_000000066D_Sub0000000002(.i_data_1(A[205][2]), .i_data_2(B[205][2]), .o_data(mult_result_r[205][2]), .i_clk(i_clk));
Sub0000000002  u_000000066E_Sub0000000002(.i_data_1(B[205][2]), .i_data_2(C[205][2]), .o_data(mult_result_i[205][2]), .i_clk(i_clk));
Sub0000000002  u_000000066F_Sub0000000002(.i_data_1(A[205][3]), .i_data_2(B[205][3]), .o_data(mult_result_r[205][3]), .i_clk(i_clk));
Sub0000000002  u_0000000670_Sub0000000002(.i_data_1(B[205][3]), .i_data_2(C[205][3]), .o_data(mult_result_i[205][3]), .i_clk(i_clk));
Sub0000000002  u_0000000671_Sub0000000002(.i_data_1(A[206][0]), .i_data_2(B[206][0]), .o_data(mult_result_r[206][0]), .i_clk(i_clk));
Sub0000000002  u_0000000672_Sub0000000002(.i_data_1(B[206][0]), .i_data_2(C[206][0]), .o_data(mult_result_i[206][0]), .i_clk(i_clk));
Sub0000000002  u_0000000673_Sub0000000002(.i_data_1(A[206][1]), .i_data_2(B[206][1]), .o_data(mult_result_r[206][1]), .i_clk(i_clk));
Sub0000000002  u_0000000674_Sub0000000002(.i_data_1(B[206][1]), .i_data_2(C[206][1]), .o_data(mult_result_i[206][1]), .i_clk(i_clk));
Sub0000000002  u_0000000675_Sub0000000002(.i_data_1(A[206][2]), .i_data_2(B[206][2]), .o_data(mult_result_r[206][2]), .i_clk(i_clk));
Sub0000000002  u_0000000676_Sub0000000002(.i_data_1(B[206][2]), .i_data_2(C[206][2]), .o_data(mult_result_i[206][2]), .i_clk(i_clk));
Sub0000000002  u_0000000677_Sub0000000002(.i_data_1(A[206][3]), .i_data_2(B[206][3]), .o_data(mult_result_r[206][3]), .i_clk(i_clk));
Sub0000000002  u_0000000678_Sub0000000002(.i_data_1(B[206][3]), .i_data_2(C[206][3]), .o_data(mult_result_i[206][3]), .i_clk(i_clk));
Sub0000000002  u_0000000679_Sub0000000002(.i_data_1(A[207][0]), .i_data_2(B[207][0]), .o_data(mult_result_r[207][0]), .i_clk(i_clk));
Sub0000000002  u_000000067A_Sub0000000002(.i_data_1(B[207][0]), .i_data_2(C[207][0]), .o_data(mult_result_i[207][0]), .i_clk(i_clk));
Sub0000000002  u_000000067B_Sub0000000002(.i_data_1(A[207][1]), .i_data_2(B[207][1]), .o_data(mult_result_r[207][1]), .i_clk(i_clk));
Sub0000000002  u_000000067C_Sub0000000002(.i_data_1(B[207][1]), .i_data_2(C[207][1]), .o_data(mult_result_i[207][1]), .i_clk(i_clk));
Sub0000000002  u_000000067D_Sub0000000002(.i_data_1(A[207][2]), .i_data_2(B[207][2]), .o_data(mult_result_r[207][2]), .i_clk(i_clk));
Sub0000000002  u_000000067E_Sub0000000002(.i_data_1(B[207][2]), .i_data_2(C[207][2]), .o_data(mult_result_i[207][2]), .i_clk(i_clk));
Sub0000000002  u_000000067F_Sub0000000002(.i_data_1(A[207][3]), .i_data_2(B[207][3]), .o_data(mult_result_r[207][3]), .i_clk(i_clk));
Sub0000000002  u_0000000680_Sub0000000002(.i_data_1(B[207][3]), .i_data_2(C[207][3]), .o_data(mult_result_i[207][3]), .i_clk(i_clk));
Sub0000000002  u_0000000681_Sub0000000002(.i_data_1(A[208][0]), .i_data_2(B[208][0]), .o_data(mult_result_r[208][0]), .i_clk(i_clk));
Sub0000000002  u_0000000682_Sub0000000002(.i_data_1(B[208][0]), .i_data_2(C[208][0]), .o_data(mult_result_i[208][0]), .i_clk(i_clk));
Sub0000000002  u_0000000683_Sub0000000002(.i_data_1(A[208][1]), .i_data_2(B[208][1]), .o_data(mult_result_r[208][1]), .i_clk(i_clk));
Sub0000000002  u_0000000684_Sub0000000002(.i_data_1(B[208][1]), .i_data_2(C[208][1]), .o_data(mult_result_i[208][1]), .i_clk(i_clk));
Sub0000000002  u_0000000685_Sub0000000002(.i_data_1(A[208][2]), .i_data_2(B[208][2]), .o_data(mult_result_r[208][2]), .i_clk(i_clk));
Sub0000000002  u_0000000686_Sub0000000002(.i_data_1(B[208][2]), .i_data_2(C[208][2]), .o_data(mult_result_i[208][2]), .i_clk(i_clk));
Sub0000000002  u_0000000687_Sub0000000002(.i_data_1(A[208][3]), .i_data_2(B[208][3]), .o_data(mult_result_r[208][3]), .i_clk(i_clk));
Sub0000000002  u_0000000688_Sub0000000002(.i_data_1(B[208][3]), .i_data_2(C[208][3]), .o_data(mult_result_i[208][3]), .i_clk(i_clk));
Sub0000000002  u_0000000689_Sub0000000002(.i_data_1(A[209][0]), .i_data_2(B[209][0]), .o_data(mult_result_r[209][0]), .i_clk(i_clk));
Sub0000000002  u_000000068A_Sub0000000002(.i_data_1(B[209][0]), .i_data_2(C[209][0]), .o_data(mult_result_i[209][0]), .i_clk(i_clk));
Sub0000000002  u_000000068B_Sub0000000002(.i_data_1(A[209][1]), .i_data_2(B[209][1]), .o_data(mult_result_r[209][1]), .i_clk(i_clk));
Sub0000000002  u_000000068C_Sub0000000002(.i_data_1(B[209][1]), .i_data_2(C[209][1]), .o_data(mult_result_i[209][1]), .i_clk(i_clk));
Sub0000000002  u_000000068D_Sub0000000002(.i_data_1(A[209][2]), .i_data_2(B[209][2]), .o_data(mult_result_r[209][2]), .i_clk(i_clk));
Sub0000000002  u_000000068E_Sub0000000002(.i_data_1(B[209][2]), .i_data_2(C[209][2]), .o_data(mult_result_i[209][2]), .i_clk(i_clk));
Sub0000000002  u_000000068F_Sub0000000002(.i_data_1(A[209][3]), .i_data_2(B[209][3]), .o_data(mult_result_r[209][3]), .i_clk(i_clk));
Sub0000000002  u_0000000690_Sub0000000002(.i_data_1(B[209][3]), .i_data_2(C[209][3]), .o_data(mult_result_i[209][3]), .i_clk(i_clk));
Sub0000000002  u_0000000691_Sub0000000002(.i_data_1(A[210][0]), .i_data_2(B[210][0]), .o_data(mult_result_r[210][0]), .i_clk(i_clk));
Sub0000000002  u_0000000692_Sub0000000002(.i_data_1(B[210][0]), .i_data_2(C[210][0]), .o_data(mult_result_i[210][0]), .i_clk(i_clk));
Sub0000000002  u_0000000693_Sub0000000002(.i_data_1(A[210][1]), .i_data_2(B[210][1]), .o_data(mult_result_r[210][1]), .i_clk(i_clk));
Sub0000000002  u_0000000694_Sub0000000002(.i_data_1(B[210][1]), .i_data_2(C[210][1]), .o_data(mult_result_i[210][1]), .i_clk(i_clk));
Sub0000000002  u_0000000695_Sub0000000002(.i_data_1(A[210][2]), .i_data_2(B[210][2]), .o_data(mult_result_r[210][2]), .i_clk(i_clk));
Sub0000000002  u_0000000696_Sub0000000002(.i_data_1(B[210][2]), .i_data_2(C[210][2]), .o_data(mult_result_i[210][2]), .i_clk(i_clk));
Sub0000000002  u_0000000697_Sub0000000002(.i_data_1(A[210][3]), .i_data_2(B[210][3]), .o_data(mult_result_r[210][3]), .i_clk(i_clk));
Sub0000000002  u_0000000698_Sub0000000002(.i_data_1(B[210][3]), .i_data_2(C[210][3]), .o_data(mult_result_i[210][3]), .i_clk(i_clk));
Sub0000000002  u_0000000699_Sub0000000002(.i_data_1(A[211][0]), .i_data_2(B[211][0]), .o_data(mult_result_r[211][0]), .i_clk(i_clk));
Sub0000000002  u_000000069A_Sub0000000002(.i_data_1(B[211][0]), .i_data_2(C[211][0]), .o_data(mult_result_i[211][0]), .i_clk(i_clk));
Sub0000000002  u_000000069B_Sub0000000002(.i_data_1(A[211][1]), .i_data_2(B[211][1]), .o_data(mult_result_r[211][1]), .i_clk(i_clk));
Sub0000000002  u_000000069C_Sub0000000002(.i_data_1(B[211][1]), .i_data_2(C[211][1]), .o_data(mult_result_i[211][1]), .i_clk(i_clk));
Sub0000000002  u_000000069D_Sub0000000002(.i_data_1(A[211][2]), .i_data_2(B[211][2]), .o_data(mult_result_r[211][2]), .i_clk(i_clk));
Sub0000000002  u_000000069E_Sub0000000002(.i_data_1(B[211][2]), .i_data_2(C[211][2]), .o_data(mult_result_i[211][2]), .i_clk(i_clk));
Sub0000000002  u_000000069F_Sub0000000002(.i_data_1(A[211][3]), .i_data_2(B[211][3]), .o_data(mult_result_r[211][3]), .i_clk(i_clk));
Sub0000000002  u_00000006A0_Sub0000000002(.i_data_1(B[211][3]), .i_data_2(C[211][3]), .o_data(mult_result_i[211][3]), .i_clk(i_clk));
Sub0000000002  u_00000006A1_Sub0000000002(.i_data_1(A[212][0]), .i_data_2(B[212][0]), .o_data(mult_result_r[212][0]), .i_clk(i_clk));
Sub0000000002  u_00000006A2_Sub0000000002(.i_data_1(B[212][0]), .i_data_2(C[212][0]), .o_data(mult_result_i[212][0]), .i_clk(i_clk));
Sub0000000002  u_00000006A3_Sub0000000002(.i_data_1(A[212][1]), .i_data_2(B[212][1]), .o_data(mult_result_r[212][1]), .i_clk(i_clk));
Sub0000000002  u_00000006A4_Sub0000000002(.i_data_1(B[212][1]), .i_data_2(C[212][1]), .o_data(mult_result_i[212][1]), .i_clk(i_clk));
Sub0000000002  u_00000006A5_Sub0000000002(.i_data_1(A[212][2]), .i_data_2(B[212][2]), .o_data(mult_result_r[212][2]), .i_clk(i_clk));
Sub0000000002  u_00000006A6_Sub0000000002(.i_data_1(B[212][2]), .i_data_2(C[212][2]), .o_data(mult_result_i[212][2]), .i_clk(i_clk));
Sub0000000002  u_00000006A7_Sub0000000002(.i_data_1(A[212][3]), .i_data_2(B[212][3]), .o_data(mult_result_r[212][3]), .i_clk(i_clk));
Sub0000000002  u_00000006A8_Sub0000000002(.i_data_1(B[212][3]), .i_data_2(C[212][3]), .o_data(mult_result_i[212][3]), .i_clk(i_clk));
Sub0000000002  u_00000006A9_Sub0000000002(.i_data_1(A[213][0]), .i_data_2(B[213][0]), .o_data(mult_result_r[213][0]), .i_clk(i_clk));
Sub0000000002  u_00000006AA_Sub0000000002(.i_data_1(B[213][0]), .i_data_2(C[213][0]), .o_data(mult_result_i[213][0]), .i_clk(i_clk));
Sub0000000002  u_00000006AB_Sub0000000002(.i_data_1(A[213][1]), .i_data_2(B[213][1]), .o_data(mult_result_r[213][1]), .i_clk(i_clk));
Sub0000000002  u_00000006AC_Sub0000000002(.i_data_1(B[213][1]), .i_data_2(C[213][1]), .o_data(mult_result_i[213][1]), .i_clk(i_clk));
Sub0000000002  u_00000006AD_Sub0000000002(.i_data_1(A[213][2]), .i_data_2(B[213][2]), .o_data(mult_result_r[213][2]), .i_clk(i_clk));
Sub0000000002  u_00000006AE_Sub0000000002(.i_data_1(B[213][2]), .i_data_2(C[213][2]), .o_data(mult_result_i[213][2]), .i_clk(i_clk));
Sub0000000002  u_00000006AF_Sub0000000002(.i_data_1(A[213][3]), .i_data_2(B[213][3]), .o_data(mult_result_r[213][3]), .i_clk(i_clk));
Sub0000000002  u_00000006B0_Sub0000000002(.i_data_1(B[213][3]), .i_data_2(C[213][3]), .o_data(mult_result_i[213][3]), .i_clk(i_clk));
Sub0000000002  u_00000006B1_Sub0000000002(.i_data_1(A[214][0]), .i_data_2(B[214][0]), .o_data(mult_result_r[214][0]), .i_clk(i_clk));
Sub0000000002  u_00000006B2_Sub0000000002(.i_data_1(B[214][0]), .i_data_2(C[214][0]), .o_data(mult_result_i[214][0]), .i_clk(i_clk));
Sub0000000002  u_00000006B3_Sub0000000002(.i_data_1(A[214][1]), .i_data_2(B[214][1]), .o_data(mult_result_r[214][1]), .i_clk(i_clk));
Sub0000000002  u_00000006B4_Sub0000000002(.i_data_1(B[214][1]), .i_data_2(C[214][1]), .o_data(mult_result_i[214][1]), .i_clk(i_clk));
Sub0000000002  u_00000006B5_Sub0000000002(.i_data_1(A[214][2]), .i_data_2(B[214][2]), .o_data(mult_result_r[214][2]), .i_clk(i_clk));
Sub0000000002  u_00000006B6_Sub0000000002(.i_data_1(B[214][2]), .i_data_2(C[214][2]), .o_data(mult_result_i[214][2]), .i_clk(i_clk));
Sub0000000002  u_00000006B7_Sub0000000002(.i_data_1(A[214][3]), .i_data_2(B[214][3]), .o_data(mult_result_r[214][3]), .i_clk(i_clk));
Sub0000000002  u_00000006B8_Sub0000000002(.i_data_1(B[214][3]), .i_data_2(C[214][3]), .o_data(mult_result_i[214][3]), .i_clk(i_clk));
Sub0000000002  u_00000006B9_Sub0000000002(.i_data_1(A[215][0]), .i_data_2(B[215][0]), .o_data(mult_result_r[215][0]), .i_clk(i_clk));
Sub0000000002  u_00000006BA_Sub0000000002(.i_data_1(B[215][0]), .i_data_2(C[215][0]), .o_data(mult_result_i[215][0]), .i_clk(i_clk));
Sub0000000002  u_00000006BB_Sub0000000002(.i_data_1(A[215][1]), .i_data_2(B[215][1]), .o_data(mult_result_r[215][1]), .i_clk(i_clk));
Sub0000000002  u_00000006BC_Sub0000000002(.i_data_1(B[215][1]), .i_data_2(C[215][1]), .o_data(mult_result_i[215][1]), .i_clk(i_clk));
Sub0000000002  u_00000006BD_Sub0000000002(.i_data_1(A[215][2]), .i_data_2(B[215][2]), .o_data(mult_result_r[215][2]), .i_clk(i_clk));
Sub0000000002  u_00000006BE_Sub0000000002(.i_data_1(B[215][2]), .i_data_2(C[215][2]), .o_data(mult_result_i[215][2]), .i_clk(i_clk));
Sub0000000002  u_00000006BF_Sub0000000002(.i_data_1(A[215][3]), .i_data_2(B[215][3]), .o_data(mult_result_r[215][3]), .i_clk(i_clk));
Sub0000000002  u_00000006C0_Sub0000000002(.i_data_1(B[215][3]), .i_data_2(C[215][3]), .o_data(mult_result_i[215][3]), .i_clk(i_clk));
Sub0000000002  u_00000006C1_Sub0000000002(.i_data_1(A[216][0]), .i_data_2(B[216][0]), .o_data(mult_result_r[216][0]), .i_clk(i_clk));
Sub0000000002  u_00000006C2_Sub0000000002(.i_data_1(B[216][0]), .i_data_2(C[216][0]), .o_data(mult_result_i[216][0]), .i_clk(i_clk));
Sub0000000002  u_00000006C3_Sub0000000002(.i_data_1(A[216][1]), .i_data_2(B[216][1]), .o_data(mult_result_r[216][1]), .i_clk(i_clk));
Sub0000000002  u_00000006C4_Sub0000000002(.i_data_1(B[216][1]), .i_data_2(C[216][1]), .o_data(mult_result_i[216][1]), .i_clk(i_clk));
Sub0000000002  u_00000006C5_Sub0000000002(.i_data_1(A[216][2]), .i_data_2(B[216][2]), .o_data(mult_result_r[216][2]), .i_clk(i_clk));
Sub0000000002  u_00000006C6_Sub0000000002(.i_data_1(B[216][2]), .i_data_2(C[216][2]), .o_data(mult_result_i[216][2]), .i_clk(i_clk));
Sub0000000002  u_00000006C7_Sub0000000002(.i_data_1(A[216][3]), .i_data_2(B[216][3]), .o_data(mult_result_r[216][3]), .i_clk(i_clk));
Sub0000000002  u_00000006C8_Sub0000000002(.i_data_1(B[216][3]), .i_data_2(C[216][3]), .o_data(mult_result_i[216][3]), .i_clk(i_clk));
Sub0000000002  u_00000006C9_Sub0000000002(.i_data_1(A[217][0]), .i_data_2(B[217][0]), .o_data(mult_result_r[217][0]), .i_clk(i_clk));
Sub0000000002  u_00000006CA_Sub0000000002(.i_data_1(B[217][0]), .i_data_2(C[217][0]), .o_data(mult_result_i[217][0]), .i_clk(i_clk));
Sub0000000002  u_00000006CB_Sub0000000002(.i_data_1(A[217][1]), .i_data_2(B[217][1]), .o_data(mult_result_r[217][1]), .i_clk(i_clk));
Sub0000000002  u_00000006CC_Sub0000000002(.i_data_1(B[217][1]), .i_data_2(C[217][1]), .o_data(mult_result_i[217][1]), .i_clk(i_clk));
Sub0000000002  u_00000006CD_Sub0000000002(.i_data_1(A[217][2]), .i_data_2(B[217][2]), .o_data(mult_result_r[217][2]), .i_clk(i_clk));
Sub0000000002  u_00000006CE_Sub0000000002(.i_data_1(B[217][2]), .i_data_2(C[217][2]), .o_data(mult_result_i[217][2]), .i_clk(i_clk));
Sub0000000002  u_00000006CF_Sub0000000002(.i_data_1(A[217][3]), .i_data_2(B[217][3]), .o_data(mult_result_r[217][3]), .i_clk(i_clk));
Sub0000000002  u_00000006D0_Sub0000000002(.i_data_1(B[217][3]), .i_data_2(C[217][3]), .o_data(mult_result_i[217][3]), .i_clk(i_clk));
Sub0000000002  u_00000006D1_Sub0000000002(.i_data_1(A[218][0]), .i_data_2(B[218][0]), .o_data(mult_result_r[218][0]), .i_clk(i_clk));
Sub0000000002  u_00000006D2_Sub0000000002(.i_data_1(B[218][0]), .i_data_2(C[218][0]), .o_data(mult_result_i[218][0]), .i_clk(i_clk));
Sub0000000002  u_00000006D3_Sub0000000002(.i_data_1(A[218][1]), .i_data_2(B[218][1]), .o_data(mult_result_r[218][1]), .i_clk(i_clk));
Sub0000000002  u_00000006D4_Sub0000000002(.i_data_1(B[218][1]), .i_data_2(C[218][1]), .o_data(mult_result_i[218][1]), .i_clk(i_clk));
Sub0000000002  u_00000006D5_Sub0000000002(.i_data_1(A[218][2]), .i_data_2(B[218][2]), .o_data(mult_result_r[218][2]), .i_clk(i_clk));
Sub0000000002  u_00000006D6_Sub0000000002(.i_data_1(B[218][2]), .i_data_2(C[218][2]), .o_data(mult_result_i[218][2]), .i_clk(i_clk));
Sub0000000002  u_00000006D7_Sub0000000002(.i_data_1(A[218][3]), .i_data_2(B[218][3]), .o_data(mult_result_r[218][3]), .i_clk(i_clk));
Sub0000000002  u_00000006D8_Sub0000000002(.i_data_1(B[218][3]), .i_data_2(C[218][3]), .o_data(mult_result_i[218][3]), .i_clk(i_clk));
Sub0000000002  u_00000006D9_Sub0000000002(.i_data_1(A[219][0]), .i_data_2(B[219][0]), .o_data(mult_result_r[219][0]), .i_clk(i_clk));
Sub0000000002  u_00000006DA_Sub0000000002(.i_data_1(B[219][0]), .i_data_2(C[219][0]), .o_data(mult_result_i[219][0]), .i_clk(i_clk));
Sub0000000002  u_00000006DB_Sub0000000002(.i_data_1(A[219][1]), .i_data_2(B[219][1]), .o_data(mult_result_r[219][1]), .i_clk(i_clk));
Sub0000000002  u_00000006DC_Sub0000000002(.i_data_1(B[219][1]), .i_data_2(C[219][1]), .o_data(mult_result_i[219][1]), .i_clk(i_clk));
Sub0000000002  u_00000006DD_Sub0000000002(.i_data_1(A[219][2]), .i_data_2(B[219][2]), .o_data(mult_result_r[219][2]), .i_clk(i_clk));
Sub0000000002  u_00000006DE_Sub0000000002(.i_data_1(B[219][2]), .i_data_2(C[219][2]), .o_data(mult_result_i[219][2]), .i_clk(i_clk));
Sub0000000002  u_00000006DF_Sub0000000002(.i_data_1(A[219][3]), .i_data_2(B[219][3]), .o_data(mult_result_r[219][3]), .i_clk(i_clk));
Sub0000000002  u_00000006E0_Sub0000000002(.i_data_1(B[219][3]), .i_data_2(C[219][3]), .o_data(mult_result_i[219][3]), .i_clk(i_clk));
Sub0000000002  u_00000006E1_Sub0000000002(.i_data_1(A[220][0]), .i_data_2(B[220][0]), .o_data(mult_result_r[220][0]), .i_clk(i_clk));
Sub0000000002  u_00000006E2_Sub0000000002(.i_data_1(B[220][0]), .i_data_2(C[220][0]), .o_data(mult_result_i[220][0]), .i_clk(i_clk));
Sub0000000002  u_00000006E3_Sub0000000002(.i_data_1(A[220][1]), .i_data_2(B[220][1]), .o_data(mult_result_r[220][1]), .i_clk(i_clk));
Sub0000000002  u_00000006E4_Sub0000000002(.i_data_1(B[220][1]), .i_data_2(C[220][1]), .o_data(mult_result_i[220][1]), .i_clk(i_clk));
Sub0000000002  u_00000006E5_Sub0000000002(.i_data_1(A[220][2]), .i_data_2(B[220][2]), .o_data(mult_result_r[220][2]), .i_clk(i_clk));
Sub0000000002  u_00000006E6_Sub0000000002(.i_data_1(B[220][2]), .i_data_2(C[220][2]), .o_data(mult_result_i[220][2]), .i_clk(i_clk));
Sub0000000002  u_00000006E7_Sub0000000002(.i_data_1(A[220][3]), .i_data_2(B[220][3]), .o_data(mult_result_r[220][3]), .i_clk(i_clk));
Sub0000000002  u_00000006E8_Sub0000000002(.i_data_1(B[220][3]), .i_data_2(C[220][3]), .o_data(mult_result_i[220][3]), .i_clk(i_clk));
Sub0000000002  u_00000006E9_Sub0000000002(.i_data_1(A[221][0]), .i_data_2(B[221][0]), .o_data(mult_result_r[221][0]), .i_clk(i_clk));
Sub0000000002  u_00000006EA_Sub0000000002(.i_data_1(B[221][0]), .i_data_2(C[221][0]), .o_data(mult_result_i[221][0]), .i_clk(i_clk));
Sub0000000002  u_00000006EB_Sub0000000002(.i_data_1(A[221][1]), .i_data_2(B[221][1]), .o_data(mult_result_r[221][1]), .i_clk(i_clk));
Sub0000000002  u_00000006EC_Sub0000000002(.i_data_1(B[221][1]), .i_data_2(C[221][1]), .o_data(mult_result_i[221][1]), .i_clk(i_clk));
Sub0000000002  u_00000006ED_Sub0000000002(.i_data_1(A[221][2]), .i_data_2(B[221][2]), .o_data(mult_result_r[221][2]), .i_clk(i_clk));
Sub0000000002  u_00000006EE_Sub0000000002(.i_data_1(B[221][2]), .i_data_2(C[221][2]), .o_data(mult_result_i[221][2]), .i_clk(i_clk));
Sub0000000002  u_00000006EF_Sub0000000002(.i_data_1(A[221][3]), .i_data_2(B[221][3]), .o_data(mult_result_r[221][3]), .i_clk(i_clk));
Sub0000000002  u_00000006F0_Sub0000000002(.i_data_1(B[221][3]), .i_data_2(C[221][3]), .o_data(mult_result_i[221][3]), .i_clk(i_clk));
Sub0000000002  u_00000006F1_Sub0000000002(.i_data_1(A[222][0]), .i_data_2(B[222][0]), .o_data(mult_result_r[222][0]), .i_clk(i_clk));
Sub0000000002  u_00000006F2_Sub0000000002(.i_data_1(B[222][0]), .i_data_2(C[222][0]), .o_data(mult_result_i[222][0]), .i_clk(i_clk));
Sub0000000002  u_00000006F3_Sub0000000002(.i_data_1(A[222][1]), .i_data_2(B[222][1]), .o_data(mult_result_r[222][1]), .i_clk(i_clk));
Sub0000000002  u_00000006F4_Sub0000000002(.i_data_1(B[222][1]), .i_data_2(C[222][1]), .o_data(mult_result_i[222][1]), .i_clk(i_clk));
Sub0000000002  u_00000006F5_Sub0000000002(.i_data_1(A[222][2]), .i_data_2(B[222][2]), .o_data(mult_result_r[222][2]), .i_clk(i_clk));
Sub0000000002  u_00000006F6_Sub0000000002(.i_data_1(B[222][2]), .i_data_2(C[222][2]), .o_data(mult_result_i[222][2]), .i_clk(i_clk));
Sub0000000002  u_00000006F7_Sub0000000002(.i_data_1(A[222][3]), .i_data_2(B[222][3]), .o_data(mult_result_r[222][3]), .i_clk(i_clk));
Sub0000000002  u_00000006F8_Sub0000000002(.i_data_1(B[222][3]), .i_data_2(C[222][3]), .o_data(mult_result_i[222][3]), .i_clk(i_clk));
Sub0000000002  u_00000006F9_Sub0000000002(.i_data_1(A[223][0]), .i_data_2(B[223][0]), .o_data(mult_result_r[223][0]), .i_clk(i_clk));
Sub0000000002  u_00000006FA_Sub0000000002(.i_data_1(B[223][0]), .i_data_2(C[223][0]), .o_data(mult_result_i[223][0]), .i_clk(i_clk));
Sub0000000002  u_00000006FB_Sub0000000002(.i_data_1(A[223][1]), .i_data_2(B[223][1]), .o_data(mult_result_r[223][1]), .i_clk(i_clk));
Sub0000000002  u_00000006FC_Sub0000000002(.i_data_1(B[223][1]), .i_data_2(C[223][1]), .o_data(mult_result_i[223][1]), .i_clk(i_clk));
Sub0000000002  u_00000006FD_Sub0000000002(.i_data_1(A[223][2]), .i_data_2(B[223][2]), .o_data(mult_result_r[223][2]), .i_clk(i_clk));
Sub0000000002  u_00000006FE_Sub0000000002(.i_data_1(B[223][2]), .i_data_2(C[223][2]), .o_data(mult_result_i[223][2]), .i_clk(i_clk));
Sub0000000002  u_00000006FF_Sub0000000002(.i_data_1(A[223][3]), .i_data_2(B[223][3]), .o_data(mult_result_r[223][3]), .i_clk(i_clk));
Sub0000000002  u_0000000700_Sub0000000002(.i_data_1(B[223][3]), .i_data_2(C[223][3]), .o_data(mult_result_i[223][3]), .i_clk(i_clk));
Sub0000000002  u_0000000701_Sub0000000002(.i_data_1(A[224][0]), .i_data_2(B[224][0]), .o_data(mult_result_r[224][0]), .i_clk(i_clk));
Sub0000000002  u_0000000702_Sub0000000002(.i_data_1(B[224][0]), .i_data_2(C[224][0]), .o_data(mult_result_i[224][0]), .i_clk(i_clk));
Sub0000000002  u_0000000703_Sub0000000002(.i_data_1(A[224][1]), .i_data_2(B[224][1]), .o_data(mult_result_r[224][1]), .i_clk(i_clk));
Sub0000000002  u_0000000704_Sub0000000002(.i_data_1(B[224][1]), .i_data_2(C[224][1]), .o_data(mult_result_i[224][1]), .i_clk(i_clk));
Sub0000000002  u_0000000705_Sub0000000002(.i_data_1(A[224][2]), .i_data_2(B[224][2]), .o_data(mult_result_r[224][2]), .i_clk(i_clk));
Sub0000000002  u_0000000706_Sub0000000002(.i_data_1(B[224][2]), .i_data_2(C[224][2]), .o_data(mult_result_i[224][2]), .i_clk(i_clk));
Sub0000000002  u_0000000707_Sub0000000002(.i_data_1(A[224][3]), .i_data_2(B[224][3]), .o_data(mult_result_r[224][3]), .i_clk(i_clk));
Sub0000000002  u_0000000708_Sub0000000002(.i_data_1(B[224][3]), .i_data_2(C[224][3]), .o_data(mult_result_i[224][3]), .i_clk(i_clk));
Sub0000000002  u_0000000709_Sub0000000002(.i_data_1(A[225][0]), .i_data_2(B[225][0]), .o_data(mult_result_r[225][0]), .i_clk(i_clk));
Sub0000000002  u_000000070A_Sub0000000002(.i_data_1(B[225][0]), .i_data_2(C[225][0]), .o_data(mult_result_i[225][0]), .i_clk(i_clk));
Sub0000000002  u_000000070B_Sub0000000002(.i_data_1(A[225][1]), .i_data_2(B[225][1]), .o_data(mult_result_r[225][1]), .i_clk(i_clk));
Sub0000000002  u_000000070C_Sub0000000002(.i_data_1(B[225][1]), .i_data_2(C[225][1]), .o_data(mult_result_i[225][1]), .i_clk(i_clk));
Sub0000000002  u_000000070D_Sub0000000002(.i_data_1(A[225][2]), .i_data_2(B[225][2]), .o_data(mult_result_r[225][2]), .i_clk(i_clk));
Sub0000000002  u_000000070E_Sub0000000002(.i_data_1(B[225][2]), .i_data_2(C[225][2]), .o_data(mult_result_i[225][2]), .i_clk(i_clk));
Sub0000000002  u_000000070F_Sub0000000002(.i_data_1(A[225][3]), .i_data_2(B[225][3]), .o_data(mult_result_r[225][3]), .i_clk(i_clk));
Sub0000000002  u_0000000710_Sub0000000002(.i_data_1(B[225][3]), .i_data_2(C[225][3]), .o_data(mult_result_i[225][3]), .i_clk(i_clk));
Sub0000000002  u_0000000711_Sub0000000002(.i_data_1(A[226][0]), .i_data_2(B[226][0]), .o_data(mult_result_r[226][0]), .i_clk(i_clk));
Sub0000000002  u_0000000712_Sub0000000002(.i_data_1(B[226][0]), .i_data_2(C[226][0]), .o_data(mult_result_i[226][0]), .i_clk(i_clk));
Sub0000000002  u_0000000713_Sub0000000002(.i_data_1(A[226][1]), .i_data_2(B[226][1]), .o_data(mult_result_r[226][1]), .i_clk(i_clk));
Sub0000000002  u_0000000714_Sub0000000002(.i_data_1(B[226][1]), .i_data_2(C[226][1]), .o_data(mult_result_i[226][1]), .i_clk(i_clk));
Sub0000000002  u_0000000715_Sub0000000002(.i_data_1(A[226][2]), .i_data_2(B[226][2]), .o_data(mult_result_r[226][2]), .i_clk(i_clk));
Sub0000000002  u_0000000716_Sub0000000002(.i_data_1(B[226][2]), .i_data_2(C[226][2]), .o_data(mult_result_i[226][2]), .i_clk(i_clk));
Sub0000000002  u_0000000717_Sub0000000002(.i_data_1(A[226][3]), .i_data_2(B[226][3]), .o_data(mult_result_r[226][3]), .i_clk(i_clk));
Sub0000000002  u_0000000718_Sub0000000002(.i_data_1(B[226][3]), .i_data_2(C[226][3]), .o_data(mult_result_i[226][3]), .i_clk(i_clk));
Sub0000000002  u_0000000719_Sub0000000002(.i_data_1(A[227][0]), .i_data_2(B[227][0]), .o_data(mult_result_r[227][0]), .i_clk(i_clk));
Sub0000000002  u_000000071A_Sub0000000002(.i_data_1(B[227][0]), .i_data_2(C[227][0]), .o_data(mult_result_i[227][0]), .i_clk(i_clk));
Sub0000000002  u_000000071B_Sub0000000002(.i_data_1(A[227][1]), .i_data_2(B[227][1]), .o_data(mult_result_r[227][1]), .i_clk(i_clk));
Sub0000000002  u_000000071C_Sub0000000002(.i_data_1(B[227][1]), .i_data_2(C[227][1]), .o_data(mult_result_i[227][1]), .i_clk(i_clk));
Sub0000000002  u_000000071D_Sub0000000002(.i_data_1(A[227][2]), .i_data_2(B[227][2]), .o_data(mult_result_r[227][2]), .i_clk(i_clk));
Sub0000000002  u_000000071E_Sub0000000002(.i_data_1(B[227][2]), .i_data_2(C[227][2]), .o_data(mult_result_i[227][2]), .i_clk(i_clk));
Sub0000000002  u_000000071F_Sub0000000002(.i_data_1(A[227][3]), .i_data_2(B[227][3]), .o_data(mult_result_r[227][3]), .i_clk(i_clk));
Sub0000000002  u_0000000720_Sub0000000002(.i_data_1(B[227][3]), .i_data_2(C[227][3]), .o_data(mult_result_i[227][3]), .i_clk(i_clk));
Sub0000000002  u_0000000721_Sub0000000002(.i_data_1(A[228][0]), .i_data_2(B[228][0]), .o_data(mult_result_r[228][0]), .i_clk(i_clk));
Sub0000000002  u_0000000722_Sub0000000002(.i_data_1(B[228][0]), .i_data_2(C[228][0]), .o_data(mult_result_i[228][0]), .i_clk(i_clk));
Sub0000000002  u_0000000723_Sub0000000002(.i_data_1(A[228][1]), .i_data_2(B[228][1]), .o_data(mult_result_r[228][1]), .i_clk(i_clk));
Sub0000000002  u_0000000724_Sub0000000002(.i_data_1(B[228][1]), .i_data_2(C[228][1]), .o_data(mult_result_i[228][1]), .i_clk(i_clk));
Sub0000000002  u_0000000725_Sub0000000002(.i_data_1(A[228][2]), .i_data_2(B[228][2]), .o_data(mult_result_r[228][2]), .i_clk(i_clk));
Sub0000000002  u_0000000726_Sub0000000002(.i_data_1(B[228][2]), .i_data_2(C[228][2]), .o_data(mult_result_i[228][2]), .i_clk(i_clk));
Sub0000000002  u_0000000727_Sub0000000002(.i_data_1(A[228][3]), .i_data_2(B[228][3]), .o_data(mult_result_r[228][3]), .i_clk(i_clk));
Sub0000000002  u_0000000728_Sub0000000002(.i_data_1(B[228][3]), .i_data_2(C[228][3]), .o_data(mult_result_i[228][3]), .i_clk(i_clk));
Sub0000000002  u_0000000729_Sub0000000002(.i_data_1(A[229][0]), .i_data_2(B[229][0]), .o_data(mult_result_r[229][0]), .i_clk(i_clk));
Sub0000000002  u_000000072A_Sub0000000002(.i_data_1(B[229][0]), .i_data_2(C[229][0]), .o_data(mult_result_i[229][0]), .i_clk(i_clk));
Sub0000000002  u_000000072B_Sub0000000002(.i_data_1(A[229][1]), .i_data_2(B[229][1]), .o_data(mult_result_r[229][1]), .i_clk(i_clk));
Sub0000000002  u_000000072C_Sub0000000002(.i_data_1(B[229][1]), .i_data_2(C[229][1]), .o_data(mult_result_i[229][1]), .i_clk(i_clk));
Sub0000000002  u_000000072D_Sub0000000002(.i_data_1(A[229][2]), .i_data_2(B[229][2]), .o_data(mult_result_r[229][2]), .i_clk(i_clk));
Sub0000000002  u_000000072E_Sub0000000002(.i_data_1(B[229][2]), .i_data_2(C[229][2]), .o_data(mult_result_i[229][2]), .i_clk(i_clk));
Sub0000000002  u_000000072F_Sub0000000002(.i_data_1(A[229][3]), .i_data_2(B[229][3]), .o_data(mult_result_r[229][3]), .i_clk(i_clk));
Sub0000000002  u_0000000730_Sub0000000002(.i_data_1(B[229][3]), .i_data_2(C[229][3]), .o_data(mult_result_i[229][3]), .i_clk(i_clk));
Sub0000000002  u_0000000731_Sub0000000002(.i_data_1(A[230][0]), .i_data_2(B[230][0]), .o_data(mult_result_r[230][0]), .i_clk(i_clk));
Sub0000000002  u_0000000732_Sub0000000002(.i_data_1(B[230][0]), .i_data_2(C[230][0]), .o_data(mult_result_i[230][0]), .i_clk(i_clk));
Sub0000000002  u_0000000733_Sub0000000002(.i_data_1(A[230][1]), .i_data_2(B[230][1]), .o_data(mult_result_r[230][1]), .i_clk(i_clk));
Sub0000000002  u_0000000734_Sub0000000002(.i_data_1(B[230][1]), .i_data_2(C[230][1]), .o_data(mult_result_i[230][1]), .i_clk(i_clk));
Sub0000000002  u_0000000735_Sub0000000002(.i_data_1(A[230][2]), .i_data_2(B[230][2]), .o_data(mult_result_r[230][2]), .i_clk(i_clk));
Sub0000000002  u_0000000736_Sub0000000002(.i_data_1(B[230][2]), .i_data_2(C[230][2]), .o_data(mult_result_i[230][2]), .i_clk(i_clk));
Sub0000000002  u_0000000737_Sub0000000002(.i_data_1(A[230][3]), .i_data_2(B[230][3]), .o_data(mult_result_r[230][3]), .i_clk(i_clk));
Sub0000000002  u_0000000738_Sub0000000002(.i_data_1(B[230][3]), .i_data_2(C[230][3]), .o_data(mult_result_i[230][3]), .i_clk(i_clk));
Sub0000000002  u_0000000739_Sub0000000002(.i_data_1(A[231][0]), .i_data_2(B[231][0]), .o_data(mult_result_r[231][0]), .i_clk(i_clk));
Sub0000000002  u_000000073A_Sub0000000002(.i_data_1(B[231][0]), .i_data_2(C[231][0]), .o_data(mult_result_i[231][0]), .i_clk(i_clk));
Sub0000000002  u_000000073B_Sub0000000002(.i_data_1(A[231][1]), .i_data_2(B[231][1]), .o_data(mult_result_r[231][1]), .i_clk(i_clk));
Sub0000000002  u_000000073C_Sub0000000002(.i_data_1(B[231][1]), .i_data_2(C[231][1]), .o_data(mult_result_i[231][1]), .i_clk(i_clk));
Sub0000000002  u_000000073D_Sub0000000002(.i_data_1(A[231][2]), .i_data_2(B[231][2]), .o_data(mult_result_r[231][2]), .i_clk(i_clk));
Sub0000000002  u_000000073E_Sub0000000002(.i_data_1(B[231][2]), .i_data_2(C[231][2]), .o_data(mult_result_i[231][2]), .i_clk(i_clk));
Sub0000000002  u_000000073F_Sub0000000002(.i_data_1(A[231][3]), .i_data_2(B[231][3]), .o_data(mult_result_r[231][3]), .i_clk(i_clk));
Sub0000000002  u_0000000740_Sub0000000002(.i_data_1(B[231][3]), .i_data_2(C[231][3]), .o_data(mult_result_i[231][3]), .i_clk(i_clk));
Sub0000000002  u_0000000741_Sub0000000002(.i_data_1(A[232][0]), .i_data_2(B[232][0]), .o_data(mult_result_r[232][0]), .i_clk(i_clk));
Sub0000000002  u_0000000742_Sub0000000002(.i_data_1(B[232][0]), .i_data_2(C[232][0]), .o_data(mult_result_i[232][0]), .i_clk(i_clk));
Sub0000000002  u_0000000743_Sub0000000002(.i_data_1(A[232][1]), .i_data_2(B[232][1]), .o_data(mult_result_r[232][1]), .i_clk(i_clk));
Sub0000000002  u_0000000744_Sub0000000002(.i_data_1(B[232][1]), .i_data_2(C[232][1]), .o_data(mult_result_i[232][1]), .i_clk(i_clk));
Sub0000000002  u_0000000745_Sub0000000002(.i_data_1(A[232][2]), .i_data_2(B[232][2]), .o_data(mult_result_r[232][2]), .i_clk(i_clk));
Sub0000000002  u_0000000746_Sub0000000002(.i_data_1(B[232][2]), .i_data_2(C[232][2]), .o_data(mult_result_i[232][2]), .i_clk(i_clk));
Sub0000000002  u_0000000747_Sub0000000002(.i_data_1(A[232][3]), .i_data_2(B[232][3]), .o_data(mult_result_r[232][3]), .i_clk(i_clk));
Sub0000000002  u_0000000748_Sub0000000002(.i_data_1(B[232][3]), .i_data_2(C[232][3]), .o_data(mult_result_i[232][3]), .i_clk(i_clk));
Sub0000000002  u_0000000749_Sub0000000002(.i_data_1(A[233][0]), .i_data_2(B[233][0]), .o_data(mult_result_r[233][0]), .i_clk(i_clk));
Sub0000000002  u_000000074A_Sub0000000002(.i_data_1(B[233][0]), .i_data_2(C[233][0]), .o_data(mult_result_i[233][0]), .i_clk(i_clk));
Sub0000000002  u_000000074B_Sub0000000002(.i_data_1(A[233][1]), .i_data_2(B[233][1]), .o_data(mult_result_r[233][1]), .i_clk(i_clk));
Sub0000000002  u_000000074C_Sub0000000002(.i_data_1(B[233][1]), .i_data_2(C[233][1]), .o_data(mult_result_i[233][1]), .i_clk(i_clk));
Sub0000000002  u_000000074D_Sub0000000002(.i_data_1(A[233][2]), .i_data_2(B[233][2]), .o_data(mult_result_r[233][2]), .i_clk(i_clk));
Sub0000000002  u_000000074E_Sub0000000002(.i_data_1(B[233][2]), .i_data_2(C[233][2]), .o_data(mult_result_i[233][2]), .i_clk(i_clk));
Sub0000000002  u_000000074F_Sub0000000002(.i_data_1(A[233][3]), .i_data_2(B[233][3]), .o_data(mult_result_r[233][3]), .i_clk(i_clk));
Sub0000000002  u_0000000750_Sub0000000002(.i_data_1(B[233][3]), .i_data_2(C[233][3]), .o_data(mult_result_i[233][3]), .i_clk(i_clk));
Sub0000000002  u_0000000751_Sub0000000002(.i_data_1(A[234][0]), .i_data_2(B[234][0]), .o_data(mult_result_r[234][0]), .i_clk(i_clk));
Sub0000000002  u_0000000752_Sub0000000002(.i_data_1(B[234][0]), .i_data_2(C[234][0]), .o_data(mult_result_i[234][0]), .i_clk(i_clk));
Sub0000000002  u_0000000753_Sub0000000002(.i_data_1(A[234][1]), .i_data_2(B[234][1]), .o_data(mult_result_r[234][1]), .i_clk(i_clk));
Sub0000000002  u_0000000754_Sub0000000002(.i_data_1(B[234][1]), .i_data_2(C[234][1]), .o_data(mult_result_i[234][1]), .i_clk(i_clk));
Sub0000000002  u_0000000755_Sub0000000002(.i_data_1(A[234][2]), .i_data_2(B[234][2]), .o_data(mult_result_r[234][2]), .i_clk(i_clk));
Sub0000000002  u_0000000756_Sub0000000002(.i_data_1(B[234][2]), .i_data_2(C[234][2]), .o_data(mult_result_i[234][2]), .i_clk(i_clk));
Sub0000000002  u_0000000757_Sub0000000002(.i_data_1(A[234][3]), .i_data_2(B[234][3]), .o_data(mult_result_r[234][3]), .i_clk(i_clk));
Sub0000000002  u_0000000758_Sub0000000002(.i_data_1(B[234][3]), .i_data_2(C[234][3]), .o_data(mult_result_i[234][3]), .i_clk(i_clk));
Sub0000000002  u_0000000759_Sub0000000002(.i_data_1(A[235][0]), .i_data_2(B[235][0]), .o_data(mult_result_r[235][0]), .i_clk(i_clk));
Sub0000000002  u_000000075A_Sub0000000002(.i_data_1(B[235][0]), .i_data_2(C[235][0]), .o_data(mult_result_i[235][0]), .i_clk(i_clk));
Sub0000000002  u_000000075B_Sub0000000002(.i_data_1(A[235][1]), .i_data_2(B[235][1]), .o_data(mult_result_r[235][1]), .i_clk(i_clk));
Sub0000000002  u_000000075C_Sub0000000002(.i_data_1(B[235][1]), .i_data_2(C[235][1]), .o_data(mult_result_i[235][1]), .i_clk(i_clk));
Sub0000000002  u_000000075D_Sub0000000002(.i_data_1(A[235][2]), .i_data_2(B[235][2]), .o_data(mult_result_r[235][2]), .i_clk(i_clk));
Sub0000000002  u_000000075E_Sub0000000002(.i_data_1(B[235][2]), .i_data_2(C[235][2]), .o_data(mult_result_i[235][2]), .i_clk(i_clk));
Sub0000000002  u_000000075F_Sub0000000002(.i_data_1(A[235][3]), .i_data_2(B[235][3]), .o_data(mult_result_r[235][3]), .i_clk(i_clk));
Sub0000000002  u_0000000760_Sub0000000002(.i_data_1(B[235][3]), .i_data_2(C[235][3]), .o_data(mult_result_i[235][3]), .i_clk(i_clk));
Sub0000000002  u_0000000761_Sub0000000002(.i_data_1(A[236][0]), .i_data_2(B[236][0]), .o_data(mult_result_r[236][0]), .i_clk(i_clk));
Sub0000000002  u_0000000762_Sub0000000002(.i_data_1(B[236][0]), .i_data_2(C[236][0]), .o_data(mult_result_i[236][0]), .i_clk(i_clk));
Sub0000000002  u_0000000763_Sub0000000002(.i_data_1(A[236][1]), .i_data_2(B[236][1]), .o_data(mult_result_r[236][1]), .i_clk(i_clk));
Sub0000000002  u_0000000764_Sub0000000002(.i_data_1(B[236][1]), .i_data_2(C[236][1]), .o_data(mult_result_i[236][1]), .i_clk(i_clk));
Sub0000000002  u_0000000765_Sub0000000002(.i_data_1(A[236][2]), .i_data_2(B[236][2]), .o_data(mult_result_r[236][2]), .i_clk(i_clk));
Sub0000000002  u_0000000766_Sub0000000002(.i_data_1(B[236][2]), .i_data_2(C[236][2]), .o_data(mult_result_i[236][2]), .i_clk(i_clk));
Sub0000000002  u_0000000767_Sub0000000002(.i_data_1(A[236][3]), .i_data_2(B[236][3]), .o_data(mult_result_r[236][3]), .i_clk(i_clk));
Sub0000000002  u_0000000768_Sub0000000002(.i_data_1(B[236][3]), .i_data_2(C[236][3]), .o_data(mult_result_i[236][3]), .i_clk(i_clk));
Sub0000000002  u_0000000769_Sub0000000002(.i_data_1(A[237][0]), .i_data_2(B[237][0]), .o_data(mult_result_r[237][0]), .i_clk(i_clk));
Sub0000000002  u_000000076A_Sub0000000002(.i_data_1(B[237][0]), .i_data_2(C[237][0]), .o_data(mult_result_i[237][0]), .i_clk(i_clk));
Sub0000000002  u_000000076B_Sub0000000002(.i_data_1(A[237][1]), .i_data_2(B[237][1]), .o_data(mult_result_r[237][1]), .i_clk(i_clk));
Sub0000000002  u_000000076C_Sub0000000002(.i_data_1(B[237][1]), .i_data_2(C[237][1]), .o_data(mult_result_i[237][1]), .i_clk(i_clk));
Sub0000000002  u_000000076D_Sub0000000002(.i_data_1(A[237][2]), .i_data_2(B[237][2]), .o_data(mult_result_r[237][2]), .i_clk(i_clk));
Sub0000000002  u_000000076E_Sub0000000002(.i_data_1(B[237][2]), .i_data_2(C[237][2]), .o_data(mult_result_i[237][2]), .i_clk(i_clk));
Sub0000000002  u_000000076F_Sub0000000002(.i_data_1(A[237][3]), .i_data_2(B[237][3]), .o_data(mult_result_r[237][3]), .i_clk(i_clk));
Sub0000000002  u_0000000770_Sub0000000002(.i_data_1(B[237][3]), .i_data_2(C[237][3]), .o_data(mult_result_i[237][3]), .i_clk(i_clk));
Sub0000000002  u_0000000771_Sub0000000002(.i_data_1(A[238][0]), .i_data_2(B[238][0]), .o_data(mult_result_r[238][0]), .i_clk(i_clk));
Sub0000000002  u_0000000772_Sub0000000002(.i_data_1(B[238][0]), .i_data_2(C[238][0]), .o_data(mult_result_i[238][0]), .i_clk(i_clk));
Sub0000000002  u_0000000773_Sub0000000002(.i_data_1(A[238][1]), .i_data_2(B[238][1]), .o_data(mult_result_r[238][1]), .i_clk(i_clk));
Sub0000000002  u_0000000774_Sub0000000002(.i_data_1(B[238][1]), .i_data_2(C[238][1]), .o_data(mult_result_i[238][1]), .i_clk(i_clk));
Sub0000000002  u_0000000775_Sub0000000002(.i_data_1(A[238][2]), .i_data_2(B[238][2]), .o_data(mult_result_r[238][2]), .i_clk(i_clk));
Sub0000000002  u_0000000776_Sub0000000002(.i_data_1(B[238][2]), .i_data_2(C[238][2]), .o_data(mult_result_i[238][2]), .i_clk(i_clk));
Sub0000000002  u_0000000777_Sub0000000002(.i_data_1(A[238][3]), .i_data_2(B[238][3]), .o_data(mult_result_r[238][3]), .i_clk(i_clk));
Sub0000000002  u_0000000778_Sub0000000002(.i_data_1(B[238][3]), .i_data_2(C[238][3]), .o_data(mult_result_i[238][3]), .i_clk(i_clk));
Sub0000000002  u_0000000779_Sub0000000002(.i_data_1(A[239][0]), .i_data_2(B[239][0]), .o_data(mult_result_r[239][0]), .i_clk(i_clk));
Sub0000000002  u_000000077A_Sub0000000002(.i_data_1(B[239][0]), .i_data_2(C[239][0]), .o_data(mult_result_i[239][0]), .i_clk(i_clk));
Sub0000000002  u_000000077B_Sub0000000002(.i_data_1(A[239][1]), .i_data_2(B[239][1]), .o_data(mult_result_r[239][1]), .i_clk(i_clk));
Sub0000000002  u_000000077C_Sub0000000002(.i_data_1(B[239][1]), .i_data_2(C[239][1]), .o_data(mult_result_i[239][1]), .i_clk(i_clk));
Sub0000000002  u_000000077D_Sub0000000002(.i_data_1(A[239][2]), .i_data_2(B[239][2]), .o_data(mult_result_r[239][2]), .i_clk(i_clk));
Sub0000000002  u_000000077E_Sub0000000002(.i_data_1(B[239][2]), .i_data_2(C[239][2]), .o_data(mult_result_i[239][2]), .i_clk(i_clk));
Sub0000000002  u_000000077F_Sub0000000002(.i_data_1(A[239][3]), .i_data_2(B[239][3]), .o_data(mult_result_r[239][3]), .i_clk(i_clk));
Sub0000000002  u_0000000780_Sub0000000002(.i_data_1(B[239][3]), .i_data_2(C[239][3]), .o_data(mult_result_i[239][3]), .i_clk(i_clk));
Sub0000000002  u_0000000781_Sub0000000002(.i_data_1(A[240][0]), .i_data_2(B[240][0]), .o_data(mult_result_r[240][0]), .i_clk(i_clk));
Sub0000000002  u_0000000782_Sub0000000002(.i_data_1(B[240][0]), .i_data_2(C[240][0]), .o_data(mult_result_i[240][0]), .i_clk(i_clk));
Sub0000000002  u_0000000783_Sub0000000002(.i_data_1(A[240][1]), .i_data_2(B[240][1]), .o_data(mult_result_r[240][1]), .i_clk(i_clk));
Sub0000000002  u_0000000784_Sub0000000002(.i_data_1(B[240][1]), .i_data_2(C[240][1]), .o_data(mult_result_i[240][1]), .i_clk(i_clk));
Sub0000000002  u_0000000785_Sub0000000002(.i_data_1(A[240][2]), .i_data_2(B[240][2]), .o_data(mult_result_r[240][2]), .i_clk(i_clk));
Sub0000000002  u_0000000786_Sub0000000002(.i_data_1(B[240][2]), .i_data_2(C[240][2]), .o_data(mult_result_i[240][2]), .i_clk(i_clk));
Sub0000000002  u_0000000787_Sub0000000002(.i_data_1(A[240][3]), .i_data_2(B[240][3]), .o_data(mult_result_r[240][3]), .i_clk(i_clk));
Sub0000000002  u_0000000788_Sub0000000002(.i_data_1(B[240][3]), .i_data_2(C[240][3]), .o_data(mult_result_i[240][3]), .i_clk(i_clk));
Sub0000000002  u_0000000789_Sub0000000002(.i_data_1(A[241][0]), .i_data_2(B[241][0]), .o_data(mult_result_r[241][0]), .i_clk(i_clk));
Sub0000000002  u_000000078A_Sub0000000002(.i_data_1(B[241][0]), .i_data_2(C[241][0]), .o_data(mult_result_i[241][0]), .i_clk(i_clk));
Sub0000000002  u_000000078B_Sub0000000002(.i_data_1(A[241][1]), .i_data_2(B[241][1]), .o_data(mult_result_r[241][1]), .i_clk(i_clk));
Sub0000000002  u_000000078C_Sub0000000002(.i_data_1(B[241][1]), .i_data_2(C[241][1]), .o_data(mult_result_i[241][1]), .i_clk(i_clk));
Sub0000000002  u_000000078D_Sub0000000002(.i_data_1(A[241][2]), .i_data_2(B[241][2]), .o_data(mult_result_r[241][2]), .i_clk(i_clk));
Sub0000000002  u_000000078E_Sub0000000002(.i_data_1(B[241][2]), .i_data_2(C[241][2]), .o_data(mult_result_i[241][2]), .i_clk(i_clk));
Sub0000000002  u_000000078F_Sub0000000002(.i_data_1(A[241][3]), .i_data_2(B[241][3]), .o_data(mult_result_r[241][3]), .i_clk(i_clk));
Sub0000000002  u_0000000790_Sub0000000002(.i_data_1(B[241][3]), .i_data_2(C[241][3]), .o_data(mult_result_i[241][3]), .i_clk(i_clk));
Sub0000000002  u_0000000791_Sub0000000002(.i_data_1(A[242][0]), .i_data_2(B[242][0]), .o_data(mult_result_r[242][0]), .i_clk(i_clk));
Sub0000000002  u_0000000792_Sub0000000002(.i_data_1(B[242][0]), .i_data_2(C[242][0]), .o_data(mult_result_i[242][0]), .i_clk(i_clk));
Sub0000000002  u_0000000793_Sub0000000002(.i_data_1(A[242][1]), .i_data_2(B[242][1]), .o_data(mult_result_r[242][1]), .i_clk(i_clk));
Sub0000000002  u_0000000794_Sub0000000002(.i_data_1(B[242][1]), .i_data_2(C[242][1]), .o_data(mult_result_i[242][1]), .i_clk(i_clk));
Sub0000000002  u_0000000795_Sub0000000002(.i_data_1(A[242][2]), .i_data_2(B[242][2]), .o_data(mult_result_r[242][2]), .i_clk(i_clk));
Sub0000000002  u_0000000796_Sub0000000002(.i_data_1(B[242][2]), .i_data_2(C[242][2]), .o_data(mult_result_i[242][2]), .i_clk(i_clk));
Sub0000000002  u_0000000797_Sub0000000002(.i_data_1(A[242][3]), .i_data_2(B[242][3]), .o_data(mult_result_r[242][3]), .i_clk(i_clk));
Sub0000000002  u_0000000798_Sub0000000002(.i_data_1(B[242][3]), .i_data_2(C[242][3]), .o_data(mult_result_i[242][3]), .i_clk(i_clk));
Sub0000000002  u_0000000799_Sub0000000002(.i_data_1(A[243][0]), .i_data_2(B[243][0]), .o_data(mult_result_r[243][0]), .i_clk(i_clk));
Sub0000000002  u_000000079A_Sub0000000002(.i_data_1(B[243][0]), .i_data_2(C[243][0]), .o_data(mult_result_i[243][0]), .i_clk(i_clk));
Sub0000000002  u_000000079B_Sub0000000002(.i_data_1(A[243][1]), .i_data_2(B[243][1]), .o_data(mult_result_r[243][1]), .i_clk(i_clk));
Sub0000000002  u_000000079C_Sub0000000002(.i_data_1(B[243][1]), .i_data_2(C[243][1]), .o_data(mult_result_i[243][1]), .i_clk(i_clk));
Sub0000000002  u_000000079D_Sub0000000002(.i_data_1(A[243][2]), .i_data_2(B[243][2]), .o_data(mult_result_r[243][2]), .i_clk(i_clk));
Sub0000000002  u_000000079E_Sub0000000002(.i_data_1(B[243][2]), .i_data_2(C[243][2]), .o_data(mult_result_i[243][2]), .i_clk(i_clk));
Sub0000000002  u_000000079F_Sub0000000002(.i_data_1(A[243][3]), .i_data_2(B[243][3]), .o_data(mult_result_r[243][3]), .i_clk(i_clk));
Sub0000000002  u_00000007A0_Sub0000000002(.i_data_1(B[243][3]), .i_data_2(C[243][3]), .o_data(mult_result_i[243][3]), .i_clk(i_clk));
Sub0000000002  u_00000007A1_Sub0000000002(.i_data_1(A[244][0]), .i_data_2(B[244][0]), .o_data(mult_result_r[244][0]), .i_clk(i_clk));
Sub0000000002  u_00000007A2_Sub0000000002(.i_data_1(B[244][0]), .i_data_2(C[244][0]), .o_data(mult_result_i[244][0]), .i_clk(i_clk));
Sub0000000002  u_00000007A3_Sub0000000002(.i_data_1(A[244][1]), .i_data_2(B[244][1]), .o_data(mult_result_r[244][1]), .i_clk(i_clk));
Sub0000000002  u_00000007A4_Sub0000000002(.i_data_1(B[244][1]), .i_data_2(C[244][1]), .o_data(mult_result_i[244][1]), .i_clk(i_clk));
Sub0000000002  u_00000007A5_Sub0000000002(.i_data_1(A[244][2]), .i_data_2(B[244][2]), .o_data(mult_result_r[244][2]), .i_clk(i_clk));
Sub0000000002  u_00000007A6_Sub0000000002(.i_data_1(B[244][2]), .i_data_2(C[244][2]), .o_data(mult_result_i[244][2]), .i_clk(i_clk));
Sub0000000002  u_00000007A7_Sub0000000002(.i_data_1(A[244][3]), .i_data_2(B[244][3]), .o_data(mult_result_r[244][3]), .i_clk(i_clk));
Sub0000000002  u_00000007A8_Sub0000000002(.i_data_1(B[244][3]), .i_data_2(C[244][3]), .o_data(mult_result_i[244][3]), .i_clk(i_clk));
Sub0000000002  u_00000007A9_Sub0000000002(.i_data_1(A[245][0]), .i_data_2(B[245][0]), .o_data(mult_result_r[245][0]), .i_clk(i_clk));
Sub0000000002  u_00000007AA_Sub0000000002(.i_data_1(B[245][0]), .i_data_2(C[245][0]), .o_data(mult_result_i[245][0]), .i_clk(i_clk));
Sub0000000002  u_00000007AB_Sub0000000002(.i_data_1(A[245][1]), .i_data_2(B[245][1]), .o_data(mult_result_r[245][1]), .i_clk(i_clk));
Sub0000000002  u_00000007AC_Sub0000000002(.i_data_1(B[245][1]), .i_data_2(C[245][1]), .o_data(mult_result_i[245][1]), .i_clk(i_clk));
Sub0000000002  u_00000007AD_Sub0000000002(.i_data_1(A[245][2]), .i_data_2(B[245][2]), .o_data(mult_result_r[245][2]), .i_clk(i_clk));
Sub0000000002  u_00000007AE_Sub0000000002(.i_data_1(B[245][2]), .i_data_2(C[245][2]), .o_data(mult_result_i[245][2]), .i_clk(i_clk));
Sub0000000002  u_00000007AF_Sub0000000002(.i_data_1(A[245][3]), .i_data_2(B[245][3]), .o_data(mult_result_r[245][3]), .i_clk(i_clk));
Sub0000000002  u_00000007B0_Sub0000000002(.i_data_1(B[245][3]), .i_data_2(C[245][3]), .o_data(mult_result_i[245][3]), .i_clk(i_clk));
Sub0000000002  u_00000007B1_Sub0000000002(.i_data_1(A[246][0]), .i_data_2(B[246][0]), .o_data(mult_result_r[246][0]), .i_clk(i_clk));
Sub0000000002  u_00000007B2_Sub0000000002(.i_data_1(B[246][0]), .i_data_2(C[246][0]), .o_data(mult_result_i[246][0]), .i_clk(i_clk));
Sub0000000002  u_00000007B3_Sub0000000002(.i_data_1(A[246][1]), .i_data_2(B[246][1]), .o_data(mult_result_r[246][1]), .i_clk(i_clk));
Sub0000000002  u_00000007B4_Sub0000000002(.i_data_1(B[246][1]), .i_data_2(C[246][1]), .o_data(mult_result_i[246][1]), .i_clk(i_clk));
Sub0000000002  u_00000007B5_Sub0000000002(.i_data_1(A[246][2]), .i_data_2(B[246][2]), .o_data(mult_result_r[246][2]), .i_clk(i_clk));
Sub0000000002  u_00000007B6_Sub0000000002(.i_data_1(B[246][2]), .i_data_2(C[246][2]), .o_data(mult_result_i[246][2]), .i_clk(i_clk));
Sub0000000002  u_00000007B7_Sub0000000002(.i_data_1(A[246][3]), .i_data_2(B[246][3]), .o_data(mult_result_r[246][3]), .i_clk(i_clk));
Sub0000000002  u_00000007B8_Sub0000000002(.i_data_1(B[246][3]), .i_data_2(C[246][3]), .o_data(mult_result_i[246][3]), .i_clk(i_clk));
Sub0000000002  u_00000007B9_Sub0000000002(.i_data_1(A[247][0]), .i_data_2(B[247][0]), .o_data(mult_result_r[247][0]), .i_clk(i_clk));
Sub0000000002  u_00000007BA_Sub0000000002(.i_data_1(B[247][0]), .i_data_2(C[247][0]), .o_data(mult_result_i[247][0]), .i_clk(i_clk));
Sub0000000002  u_00000007BB_Sub0000000002(.i_data_1(A[247][1]), .i_data_2(B[247][1]), .o_data(mult_result_r[247][1]), .i_clk(i_clk));
Sub0000000002  u_00000007BC_Sub0000000002(.i_data_1(B[247][1]), .i_data_2(C[247][1]), .o_data(mult_result_i[247][1]), .i_clk(i_clk));
Sub0000000002  u_00000007BD_Sub0000000002(.i_data_1(A[247][2]), .i_data_2(B[247][2]), .o_data(mult_result_r[247][2]), .i_clk(i_clk));
Sub0000000002  u_00000007BE_Sub0000000002(.i_data_1(B[247][2]), .i_data_2(C[247][2]), .o_data(mult_result_i[247][2]), .i_clk(i_clk));
Sub0000000002  u_00000007BF_Sub0000000002(.i_data_1(A[247][3]), .i_data_2(B[247][3]), .o_data(mult_result_r[247][3]), .i_clk(i_clk));
Sub0000000002  u_00000007C0_Sub0000000002(.i_data_1(B[247][3]), .i_data_2(C[247][3]), .o_data(mult_result_i[247][3]), .i_clk(i_clk));
Sub0000000002  u_00000007C1_Sub0000000002(.i_data_1(A[248][0]), .i_data_2(B[248][0]), .o_data(mult_result_r[248][0]), .i_clk(i_clk));
Sub0000000002  u_00000007C2_Sub0000000002(.i_data_1(B[248][0]), .i_data_2(C[248][0]), .o_data(mult_result_i[248][0]), .i_clk(i_clk));
Sub0000000002  u_00000007C3_Sub0000000002(.i_data_1(A[248][1]), .i_data_2(B[248][1]), .o_data(mult_result_r[248][1]), .i_clk(i_clk));
Sub0000000002  u_00000007C4_Sub0000000002(.i_data_1(B[248][1]), .i_data_2(C[248][1]), .o_data(mult_result_i[248][1]), .i_clk(i_clk));
Sub0000000002  u_00000007C5_Sub0000000002(.i_data_1(A[248][2]), .i_data_2(B[248][2]), .o_data(mult_result_r[248][2]), .i_clk(i_clk));
Sub0000000002  u_00000007C6_Sub0000000002(.i_data_1(B[248][2]), .i_data_2(C[248][2]), .o_data(mult_result_i[248][2]), .i_clk(i_clk));
Sub0000000002  u_00000007C7_Sub0000000002(.i_data_1(A[248][3]), .i_data_2(B[248][3]), .o_data(mult_result_r[248][3]), .i_clk(i_clk));
Sub0000000002  u_00000007C8_Sub0000000002(.i_data_1(B[248][3]), .i_data_2(C[248][3]), .o_data(mult_result_i[248][3]), .i_clk(i_clk));
Sub0000000002  u_00000007C9_Sub0000000002(.i_data_1(A[249][0]), .i_data_2(B[249][0]), .o_data(mult_result_r[249][0]), .i_clk(i_clk));
Sub0000000002  u_00000007CA_Sub0000000002(.i_data_1(B[249][0]), .i_data_2(C[249][0]), .o_data(mult_result_i[249][0]), .i_clk(i_clk));
Sub0000000002  u_00000007CB_Sub0000000002(.i_data_1(A[249][1]), .i_data_2(B[249][1]), .o_data(mult_result_r[249][1]), .i_clk(i_clk));
Sub0000000002  u_00000007CC_Sub0000000002(.i_data_1(B[249][1]), .i_data_2(C[249][1]), .o_data(mult_result_i[249][1]), .i_clk(i_clk));
Sub0000000002  u_00000007CD_Sub0000000002(.i_data_1(A[249][2]), .i_data_2(B[249][2]), .o_data(mult_result_r[249][2]), .i_clk(i_clk));
Sub0000000002  u_00000007CE_Sub0000000002(.i_data_1(B[249][2]), .i_data_2(C[249][2]), .o_data(mult_result_i[249][2]), .i_clk(i_clk));
Sub0000000002  u_00000007CF_Sub0000000002(.i_data_1(A[249][3]), .i_data_2(B[249][3]), .o_data(mult_result_r[249][3]), .i_clk(i_clk));
Sub0000000002  u_00000007D0_Sub0000000002(.i_data_1(B[249][3]), .i_data_2(C[249][3]), .o_data(mult_result_i[249][3]), .i_clk(i_clk));
Sub0000000002  u_00000007D1_Sub0000000002(.i_data_1(A[250][0]), .i_data_2(B[250][0]), .o_data(mult_result_r[250][0]), .i_clk(i_clk));
Sub0000000002  u_00000007D2_Sub0000000002(.i_data_1(B[250][0]), .i_data_2(C[250][0]), .o_data(mult_result_i[250][0]), .i_clk(i_clk));
Sub0000000002  u_00000007D3_Sub0000000002(.i_data_1(A[250][1]), .i_data_2(B[250][1]), .o_data(mult_result_r[250][1]), .i_clk(i_clk));
Sub0000000002  u_00000007D4_Sub0000000002(.i_data_1(B[250][1]), .i_data_2(C[250][1]), .o_data(mult_result_i[250][1]), .i_clk(i_clk));
Sub0000000002  u_00000007D5_Sub0000000002(.i_data_1(A[250][2]), .i_data_2(B[250][2]), .o_data(mult_result_r[250][2]), .i_clk(i_clk));
Sub0000000002  u_00000007D6_Sub0000000002(.i_data_1(B[250][2]), .i_data_2(C[250][2]), .o_data(mult_result_i[250][2]), .i_clk(i_clk));
Sub0000000002  u_00000007D7_Sub0000000002(.i_data_1(A[250][3]), .i_data_2(B[250][3]), .o_data(mult_result_r[250][3]), .i_clk(i_clk));
Sub0000000002  u_00000007D8_Sub0000000002(.i_data_1(B[250][3]), .i_data_2(C[250][3]), .o_data(mult_result_i[250][3]), .i_clk(i_clk));
Sub0000000002  u_00000007D9_Sub0000000002(.i_data_1(A[251][0]), .i_data_2(B[251][0]), .o_data(mult_result_r[251][0]), .i_clk(i_clk));
Sub0000000002  u_00000007DA_Sub0000000002(.i_data_1(B[251][0]), .i_data_2(C[251][0]), .o_data(mult_result_i[251][0]), .i_clk(i_clk));
Sub0000000002  u_00000007DB_Sub0000000002(.i_data_1(A[251][1]), .i_data_2(B[251][1]), .o_data(mult_result_r[251][1]), .i_clk(i_clk));
Sub0000000002  u_00000007DC_Sub0000000002(.i_data_1(B[251][1]), .i_data_2(C[251][1]), .o_data(mult_result_i[251][1]), .i_clk(i_clk));
Sub0000000002  u_00000007DD_Sub0000000002(.i_data_1(A[251][2]), .i_data_2(B[251][2]), .o_data(mult_result_r[251][2]), .i_clk(i_clk));
Sub0000000002  u_00000007DE_Sub0000000002(.i_data_1(B[251][2]), .i_data_2(C[251][2]), .o_data(mult_result_i[251][2]), .i_clk(i_clk));
Sub0000000002  u_00000007DF_Sub0000000002(.i_data_1(A[251][3]), .i_data_2(B[251][3]), .o_data(mult_result_r[251][3]), .i_clk(i_clk));
Sub0000000002  u_00000007E0_Sub0000000002(.i_data_1(B[251][3]), .i_data_2(C[251][3]), .o_data(mult_result_i[251][3]), .i_clk(i_clk));
Sub0000000002  u_00000007E1_Sub0000000002(.i_data_1(A[252][0]), .i_data_2(B[252][0]), .o_data(mult_result_r[252][0]), .i_clk(i_clk));
Sub0000000002  u_00000007E2_Sub0000000002(.i_data_1(B[252][0]), .i_data_2(C[252][0]), .o_data(mult_result_i[252][0]), .i_clk(i_clk));
Sub0000000002  u_00000007E3_Sub0000000002(.i_data_1(A[252][1]), .i_data_2(B[252][1]), .o_data(mult_result_r[252][1]), .i_clk(i_clk));
Sub0000000002  u_00000007E4_Sub0000000002(.i_data_1(B[252][1]), .i_data_2(C[252][1]), .o_data(mult_result_i[252][1]), .i_clk(i_clk));
Sub0000000002  u_00000007E5_Sub0000000002(.i_data_1(A[252][2]), .i_data_2(B[252][2]), .o_data(mult_result_r[252][2]), .i_clk(i_clk));
Sub0000000002  u_00000007E6_Sub0000000002(.i_data_1(B[252][2]), .i_data_2(C[252][2]), .o_data(mult_result_i[252][2]), .i_clk(i_clk));
Sub0000000002  u_00000007E7_Sub0000000002(.i_data_1(A[252][3]), .i_data_2(B[252][3]), .o_data(mult_result_r[252][3]), .i_clk(i_clk));
Sub0000000002  u_00000007E8_Sub0000000002(.i_data_1(B[252][3]), .i_data_2(C[252][3]), .o_data(mult_result_i[252][3]), .i_clk(i_clk));
Sub0000000002  u_00000007E9_Sub0000000002(.i_data_1(A[253][0]), .i_data_2(B[253][0]), .o_data(mult_result_r[253][0]), .i_clk(i_clk));
Sub0000000002  u_00000007EA_Sub0000000002(.i_data_1(B[253][0]), .i_data_2(C[253][0]), .o_data(mult_result_i[253][0]), .i_clk(i_clk));
Sub0000000002  u_00000007EB_Sub0000000002(.i_data_1(A[253][1]), .i_data_2(B[253][1]), .o_data(mult_result_r[253][1]), .i_clk(i_clk));
Sub0000000002  u_00000007EC_Sub0000000002(.i_data_1(B[253][1]), .i_data_2(C[253][1]), .o_data(mult_result_i[253][1]), .i_clk(i_clk));
Sub0000000002  u_00000007ED_Sub0000000002(.i_data_1(A[253][2]), .i_data_2(B[253][2]), .o_data(mult_result_r[253][2]), .i_clk(i_clk));
Sub0000000002  u_00000007EE_Sub0000000002(.i_data_1(B[253][2]), .i_data_2(C[253][2]), .o_data(mult_result_i[253][2]), .i_clk(i_clk));
Sub0000000002  u_00000007EF_Sub0000000002(.i_data_1(A[253][3]), .i_data_2(B[253][3]), .o_data(mult_result_r[253][3]), .i_clk(i_clk));
Sub0000000002  u_00000007F0_Sub0000000002(.i_data_1(B[253][3]), .i_data_2(C[253][3]), .o_data(mult_result_i[253][3]), .i_clk(i_clk));
Sub0000000002  u_00000007F1_Sub0000000002(.i_data_1(A[254][0]), .i_data_2(B[254][0]), .o_data(mult_result_r[254][0]), .i_clk(i_clk));
Sub0000000002  u_00000007F2_Sub0000000002(.i_data_1(B[254][0]), .i_data_2(C[254][0]), .o_data(mult_result_i[254][0]), .i_clk(i_clk));
Sub0000000002  u_00000007F3_Sub0000000002(.i_data_1(A[254][1]), .i_data_2(B[254][1]), .o_data(mult_result_r[254][1]), .i_clk(i_clk));
Sub0000000002  u_00000007F4_Sub0000000002(.i_data_1(B[254][1]), .i_data_2(C[254][1]), .o_data(mult_result_i[254][1]), .i_clk(i_clk));
Sub0000000002  u_00000007F5_Sub0000000002(.i_data_1(A[254][2]), .i_data_2(B[254][2]), .o_data(mult_result_r[254][2]), .i_clk(i_clk));
Sub0000000002  u_00000007F6_Sub0000000002(.i_data_1(B[254][2]), .i_data_2(C[254][2]), .o_data(mult_result_i[254][2]), .i_clk(i_clk));
Sub0000000002  u_00000007F7_Sub0000000002(.i_data_1(A[254][3]), .i_data_2(B[254][3]), .o_data(mult_result_r[254][3]), .i_clk(i_clk));
Sub0000000002  u_00000007F8_Sub0000000002(.i_data_1(B[254][3]), .i_data_2(C[254][3]), .o_data(mult_result_i[254][3]), .i_clk(i_clk));
Sub0000000002  u_00000007F9_Sub0000000002(.i_data_1(A[255][0]), .i_data_2(B[255][0]), .o_data(mult_result_r[255][0]), .i_clk(i_clk));
Sub0000000002  u_00000007FA_Sub0000000002(.i_data_1(B[255][0]), .i_data_2(C[255][0]), .o_data(mult_result_i[255][0]), .i_clk(i_clk));
Sub0000000002  u_00000007FB_Sub0000000002(.i_data_1(A[255][1]), .i_data_2(B[255][1]), .o_data(mult_result_r[255][1]), .i_clk(i_clk));
Sub0000000002  u_00000007FC_Sub0000000002(.i_data_1(B[255][1]), .i_data_2(C[255][1]), .o_data(mult_result_i[255][1]), .i_clk(i_clk));
Sub0000000002  u_00000007FD_Sub0000000002(.i_data_1(A[255][2]), .i_data_2(B[255][2]), .o_data(mult_result_r[255][2]), .i_clk(i_clk));
Sub0000000002  u_00000007FE_Sub0000000002(.i_data_1(B[255][2]), .i_data_2(C[255][2]), .o_data(mult_result_i[255][2]), .i_clk(i_clk));
Sub0000000002  u_00000007FF_Sub0000000002(.i_data_1(A[255][3]), .i_data_2(B[255][3]), .o_data(mult_result_r[255][3]), .i_clk(i_clk));
Sub0000000002  u_0000000800_Sub0000000002(.i_data_1(B[255][3]), .i_data_2(C[255][3]), .o_data(mult_result_i[255][3]), .i_clk(i_clk));
 wire [256*12-1:0] result_r;
 wire [256*12-1:0] result_i;
 assign o_result = {result_i, result_r};
AdderTree0000000001  u_0000000001_AdderTree0000000001(.i_data({mult_result_r[0][3],mult_result_r[0][2],mult_result_r[0][1],mult_result_r[0][0]}), .o_data(result_r[0*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000002_AdderTree0000000001(.i_data({mult_result_i[0][3],mult_result_i[0][2],mult_result_i[0][1],mult_result_i[0][0]}), .o_data(result_i[0*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000003_AdderTree0000000001(.i_data({mult_result_r[1][3],mult_result_r[1][2],mult_result_r[1][1],mult_result_r[1][0]}), .o_data(result_r[1*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000004_AdderTree0000000001(.i_data({mult_result_i[1][3],mult_result_i[1][2],mult_result_i[1][1],mult_result_i[1][0]}), .o_data(result_i[1*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000005_AdderTree0000000001(.i_data({mult_result_r[2][3],mult_result_r[2][2],mult_result_r[2][1],mult_result_r[2][0]}), .o_data(result_r[2*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000006_AdderTree0000000001(.i_data({mult_result_i[2][3],mult_result_i[2][2],mult_result_i[2][1],mult_result_i[2][0]}), .o_data(result_i[2*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000007_AdderTree0000000001(.i_data({mult_result_r[3][3],mult_result_r[3][2],mult_result_r[3][1],mult_result_r[3][0]}), .o_data(result_r[3*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000008_AdderTree0000000001(.i_data({mult_result_i[3][3],mult_result_i[3][2],mult_result_i[3][1],mult_result_i[3][0]}), .o_data(result_i[3*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000009_AdderTree0000000001(.i_data({mult_result_r[4][3],mult_result_r[4][2],mult_result_r[4][1],mult_result_r[4][0]}), .o_data(result_r[4*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000000A_AdderTree0000000001(.i_data({mult_result_i[4][3],mult_result_i[4][2],mult_result_i[4][1],mult_result_i[4][0]}), .o_data(result_i[4*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000000B_AdderTree0000000001(.i_data({mult_result_r[5][3],mult_result_r[5][2],mult_result_r[5][1],mult_result_r[5][0]}), .o_data(result_r[5*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000000C_AdderTree0000000001(.i_data({mult_result_i[5][3],mult_result_i[5][2],mult_result_i[5][1],mult_result_i[5][0]}), .o_data(result_i[5*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000000D_AdderTree0000000001(.i_data({mult_result_r[6][3],mult_result_r[6][2],mult_result_r[6][1],mult_result_r[6][0]}), .o_data(result_r[6*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000000E_AdderTree0000000001(.i_data({mult_result_i[6][3],mult_result_i[6][2],mult_result_i[6][1],mult_result_i[6][0]}), .o_data(result_i[6*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000000F_AdderTree0000000001(.i_data({mult_result_r[7][3],mult_result_r[7][2],mult_result_r[7][1],mult_result_r[7][0]}), .o_data(result_r[7*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000010_AdderTree0000000001(.i_data({mult_result_i[7][3],mult_result_i[7][2],mult_result_i[7][1],mult_result_i[7][0]}), .o_data(result_i[7*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000011_AdderTree0000000001(.i_data({mult_result_r[8][3],mult_result_r[8][2],mult_result_r[8][1],mult_result_r[8][0]}), .o_data(result_r[8*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000012_AdderTree0000000001(.i_data({mult_result_i[8][3],mult_result_i[8][2],mult_result_i[8][1],mult_result_i[8][0]}), .o_data(result_i[8*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000013_AdderTree0000000001(.i_data({mult_result_r[9][3],mult_result_r[9][2],mult_result_r[9][1],mult_result_r[9][0]}), .o_data(result_r[9*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000014_AdderTree0000000001(.i_data({mult_result_i[9][3],mult_result_i[9][2],mult_result_i[9][1],mult_result_i[9][0]}), .o_data(result_i[9*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000015_AdderTree0000000001(.i_data({mult_result_r[10][3],mult_result_r[10][2],mult_result_r[10][1],mult_result_r[10][0]}), .o_data(result_r[10*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000016_AdderTree0000000001(.i_data({mult_result_i[10][3],mult_result_i[10][2],mult_result_i[10][1],mult_result_i[10][0]}), .o_data(result_i[10*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000017_AdderTree0000000001(.i_data({mult_result_r[11][3],mult_result_r[11][2],mult_result_r[11][1],mult_result_r[11][0]}), .o_data(result_r[11*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000018_AdderTree0000000001(.i_data({mult_result_i[11][3],mult_result_i[11][2],mult_result_i[11][1],mult_result_i[11][0]}), .o_data(result_i[11*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000019_AdderTree0000000001(.i_data({mult_result_r[12][3],mult_result_r[12][2],mult_result_r[12][1],mult_result_r[12][0]}), .o_data(result_r[12*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000001A_AdderTree0000000001(.i_data({mult_result_i[12][3],mult_result_i[12][2],mult_result_i[12][1],mult_result_i[12][0]}), .o_data(result_i[12*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000001B_AdderTree0000000001(.i_data({mult_result_r[13][3],mult_result_r[13][2],mult_result_r[13][1],mult_result_r[13][0]}), .o_data(result_r[13*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000001C_AdderTree0000000001(.i_data({mult_result_i[13][3],mult_result_i[13][2],mult_result_i[13][1],mult_result_i[13][0]}), .o_data(result_i[13*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000001D_AdderTree0000000001(.i_data({mult_result_r[14][3],mult_result_r[14][2],mult_result_r[14][1],mult_result_r[14][0]}), .o_data(result_r[14*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000001E_AdderTree0000000001(.i_data({mult_result_i[14][3],mult_result_i[14][2],mult_result_i[14][1],mult_result_i[14][0]}), .o_data(result_i[14*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000001F_AdderTree0000000001(.i_data({mult_result_r[15][3],mult_result_r[15][2],mult_result_r[15][1],mult_result_r[15][0]}), .o_data(result_r[15*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000020_AdderTree0000000001(.i_data({mult_result_i[15][3],mult_result_i[15][2],mult_result_i[15][1],mult_result_i[15][0]}), .o_data(result_i[15*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000021_AdderTree0000000001(.i_data({mult_result_r[16][3],mult_result_r[16][2],mult_result_r[16][1],mult_result_r[16][0]}), .o_data(result_r[16*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000022_AdderTree0000000001(.i_data({mult_result_i[16][3],mult_result_i[16][2],mult_result_i[16][1],mult_result_i[16][0]}), .o_data(result_i[16*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000023_AdderTree0000000001(.i_data({mult_result_r[17][3],mult_result_r[17][2],mult_result_r[17][1],mult_result_r[17][0]}), .o_data(result_r[17*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000024_AdderTree0000000001(.i_data({mult_result_i[17][3],mult_result_i[17][2],mult_result_i[17][1],mult_result_i[17][0]}), .o_data(result_i[17*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000025_AdderTree0000000001(.i_data({mult_result_r[18][3],mult_result_r[18][2],mult_result_r[18][1],mult_result_r[18][0]}), .o_data(result_r[18*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000026_AdderTree0000000001(.i_data({mult_result_i[18][3],mult_result_i[18][2],mult_result_i[18][1],mult_result_i[18][0]}), .o_data(result_i[18*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000027_AdderTree0000000001(.i_data({mult_result_r[19][3],mult_result_r[19][2],mult_result_r[19][1],mult_result_r[19][0]}), .o_data(result_r[19*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000028_AdderTree0000000001(.i_data({mult_result_i[19][3],mult_result_i[19][2],mult_result_i[19][1],mult_result_i[19][0]}), .o_data(result_i[19*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000029_AdderTree0000000001(.i_data({mult_result_r[20][3],mult_result_r[20][2],mult_result_r[20][1],mult_result_r[20][0]}), .o_data(result_r[20*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000002A_AdderTree0000000001(.i_data({mult_result_i[20][3],mult_result_i[20][2],mult_result_i[20][1],mult_result_i[20][0]}), .o_data(result_i[20*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000002B_AdderTree0000000001(.i_data({mult_result_r[21][3],mult_result_r[21][2],mult_result_r[21][1],mult_result_r[21][0]}), .o_data(result_r[21*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000002C_AdderTree0000000001(.i_data({mult_result_i[21][3],mult_result_i[21][2],mult_result_i[21][1],mult_result_i[21][0]}), .o_data(result_i[21*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000002D_AdderTree0000000001(.i_data({mult_result_r[22][3],mult_result_r[22][2],mult_result_r[22][1],mult_result_r[22][0]}), .o_data(result_r[22*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000002E_AdderTree0000000001(.i_data({mult_result_i[22][3],mult_result_i[22][2],mult_result_i[22][1],mult_result_i[22][0]}), .o_data(result_i[22*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000002F_AdderTree0000000001(.i_data({mult_result_r[23][3],mult_result_r[23][2],mult_result_r[23][1],mult_result_r[23][0]}), .o_data(result_r[23*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000030_AdderTree0000000001(.i_data({mult_result_i[23][3],mult_result_i[23][2],mult_result_i[23][1],mult_result_i[23][0]}), .o_data(result_i[23*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000031_AdderTree0000000001(.i_data({mult_result_r[24][3],mult_result_r[24][2],mult_result_r[24][1],mult_result_r[24][0]}), .o_data(result_r[24*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000032_AdderTree0000000001(.i_data({mult_result_i[24][3],mult_result_i[24][2],mult_result_i[24][1],mult_result_i[24][0]}), .o_data(result_i[24*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000033_AdderTree0000000001(.i_data({mult_result_r[25][3],mult_result_r[25][2],mult_result_r[25][1],mult_result_r[25][0]}), .o_data(result_r[25*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000034_AdderTree0000000001(.i_data({mult_result_i[25][3],mult_result_i[25][2],mult_result_i[25][1],mult_result_i[25][0]}), .o_data(result_i[25*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000035_AdderTree0000000001(.i_data({mult_result_r[26][3],mult_result_r[26][2],mult_result_r[26][1],mult_result_r[26][0]}), .o_data(result_r[26*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000036_AdderTree0000000001(.i_data({mult_result_i[26][3],mult_result_i[26][2],mult_result_i[26][1],mult_result_i[26][0]}), .o_data(result_i[26*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000037_AdderTree0000000001(.i_data({mult_result_r[27][3],mult_result_r[27][2],mult_result_r[27][1],mult_result_r[27][0]}), .o_data(result_r[27*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000038_AdderTree0000000001(.i_data({mult_result_i[27][3],mult_result_i[27][2],mult_result_i[27][1],mult_result_i[27][0]}), .o_data(result_i[27*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000039_AdderTree0000000001(.i_data({mult_result_r[28][3],mult_result_r[28][2],mult_result_r[28][1],mult_result_r[28][0]}), .o_data(result_r[28*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000003A_AdderTree0000000001(.i_data({mult_result_i[28][3],mult_result_i[28][2],mult_result_i[28][1],mult_result_i[28][0]}), .o_data(result_i[28*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000003B_AdderTree0000000001(.i_data({mult_result_r[29][3],mult_result_r[29][2],mult_result_r[29][1],mult_result_r[29][0]}), .o_data(result_r[29*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000003C_AdderTree0000000001(.i_data({mult_result_i[29][3],mult_result_i[29][2],mult_result_i[29][1],mult_result_i[29][0]}), .o_data(result_i[29*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000003D_AdderTree0000000001(.i_data({mult_result_r[30][3],mult_result_r[30][2],mult_result_r[30][1],mult_result_r[30][0]}), .o_data(result_r[30*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000003E_AdderTree0000000001(.i_data({mult_result_i[30][3],mult_result_i[30][2],mult_result_i[30][1],mult_result_i[30][0]}), .o_data(result_i[30*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000003F_AdderTree0000000001(.i_data({mult_result_r[31][3],mult_result_r[31][2],mult_result_r[31][1],mult_result_r[31][0]}), .o_data(result_r[31*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000040_AdderTree0000000001(.i_data({mult_result_i[31][3],mult_result_i[31][2],mult_result_i[31][1],mult_result_i[31][0]}), .o_data(result_i[31*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000041_AdderTree0000000001(.i_data({mult_result_r[32][3],mult_result_r[32][2],mult_result_r[32][1],mult_result_r[32][0]}), .o_data(result_r[32*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000042_AdderTree0000000001(.i_data({mult_result_i[32][3],mult_result_i[32][2],mult_result_i[32][1],mult_result_i[32][0]}), .o_data(result_i[32*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000043_AdderTree0000000001(.i_data({mult_result_r[33][3],mult_result_r[33][2],mult_result_r[33][1],mult_result_r[33][0]}), .o_data(result_r[33*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000044_AdderTree0000000001(.i_data({mult_result_i[33][3],mult_result_i[33][2],mult_result_i[33][1],mult_result_i[33][0]}), .o_data(result_i[33*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000045_AdderTree0000000001(.i_data({mult_result_r[34][3],mult_result_r[34][2],mult_result_r[34][1],mult_result_r[34][0]}), .o_data(result_r[34*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000046_AdderTree0000000001(.i_data({mult_result_i[34][3],mult_result_i[34][2],mult_result_i[34][1],mult_result_i[34][0]}), .o_data(result_i[34*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000047_AdderTree0000000001(.i_data({mult_result_r[35][3],mult_result_r[35][2],mult_result_r[35][1],mult_result_r[35][0]}), .o_data(result_r[35*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000048_AdderTree0000000001(.i_data({mult_result_i[35][3],mult_result_i[35][2],mult_result_i[35][1],mult_result_i[35][0]}), .o_data(result_i[35*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000049_AdderTree0000000001(.i_data({mult_result_r[36][3],mult_result_r[36][2],mult_result_r[36][1],mult_result_r[36][0]}), .o_data(result_r[36*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000004A_AdderTree0000000001(.i_data({mult_result_i[36][3],mult_result_i[36][2],mult_result_i[36][1],mult_result_i[36][0]}), .o_data(result_i[36*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000004B_AdderTree0000000001(.i_data({mult_result_r[37][3],mult_result_r[37][2],mult_result_r[37][1],mult_result_r[37][0]}), .o_data(result_r[37*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000004C_AdderTree0000000001(.i_data({mult_result_i[37][3],mult_result_i[37][2],mult_result_i[37][1],mult_result_i[37][0]}), .o_data(result_i[37*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000004D_AdderTree0000000001(.i_data({mult_result_r[38][3],mult_result_r[38][2],mult_result_r[38][1],mult_result_r[38][0]}), .o_data(result_r[38*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000004E_AdderTree0000000001(.i_data({mult_result_i[38][3],mult_result_i[38][2],mult_result_i[38][1],mult_result_i[38][0]}), .o_data(result_i[38*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000004F_AdderTree0000000001(.i_data({mult_result_r[39][3],mult_result_r[39][2],mult_result_r[39][1],mult_result_r[39][0]}), .o_data(result_r[39*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000050_AdderTree0000000001(.i_data({mult_result_i[39][3],mult_result_i[39][2],mult_result_i[39][1],mult_result_i[39][0]}), .o_data(result_i[39*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000051_AdderTree0000000001(.i_data({mult_result_r[40][3],mult_result_r[40][2],mult_result_r[40][1],mult_result_r[40][0]}), .o_data(result_r[40*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000052_AdderTree0000000001(.i_data({mult_result_i[40][3],mult_result_i[40][2],mult_result_i[40][1],mult_result_i[40][0]}), .o_data(result_i[40*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000053_AdderTree0000000001(.i_data({mult_result_r[41][3],mult_result_r[41][2],mult_result_r[41][1],mult_result_r[41][0]}), .o_data(result_r[41*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000054_AdderTree0000000001(.i_data({mult_result_i[41][3],mult_result_i[41][2],mult_result_i[41][1],mult_result_i[41][0]}), .o_data(result_i[41*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000055_AdderTree0000000001(.i_data({mult_result_r[42][3],mult_result_r[42][2],mult_result_r[42][1],mult_result_r[42][0]}), .o_data(result_r[42*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000056_AdderTree0000000001(.i_data({mult_result_i[42][3],mult_result_i[42][2],mult_result_i[42][1],mult_result_i[42][0]}), .o_data(result_i[42*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000057_AdderTree0000000001(.i_data({mult_result_r[43][3],mult_result_r[43][2],mult_result_r[43][1],mult_result_r[43][0]}), .o_data(result_r[43*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000058_AdderTree0000000001(.i_data({mult_result_i[43][3],mult_result_i[43][2],mult_result_i[43][1],mult_result_i[43][0]}), .o_data(result_i[43*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000059_AdderTree0000000001(.i_data({mult_result_r[44][3],mult_result_r[44][2],mult_result_r[44][1],mult_result_r[44][0]}), .o_data(result_r[44*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000005A_AdderTree0000000001(.i_data({mult_result_i[44][3],mult_result_i[44][2],mult_result_i[44][1],mult_result_i[44][0]}), .o_data(result_i[44*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000005B_AdderTree0000000001(.i_data({mult_result_r[45][3],mult_result_r[45][2],mult_result_r[45][1],mult_result_r[45][0]}), .o_data(result_r[45*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000005C_AdderTree0000000001(.i_data({mult_result_i[45][3],mult_result_i[45][2],mult_result_i[45][1],mult_result_i[45][0]}), .o_data(result_i[45*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000005D_AdderTree0000000001(.i_data({mult_result_r[46][3],mult_result_r[46][2],mult_result_r[46][1],mult_result_r[46][0]}), .o_data(result_r[46*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000005E_AdderTree0000000001(.i_data({mult_result_i[46][3],mult_result_i[46][2],mult_result_i[46][1],mult_result_i[46][0]}), .o_data(result_i[46*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000005F_AdderTree0000000001(.i_data({mult_result_r[47][3],mult_result_r[47][2],mult_result_r[47][1],mult_result_r[47][0]}), .o_data(result_r[47*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000060_AdderTree0000000001(.i_data({mult_result_i[47][3],mult_result_i[47][2],mult_result_i[47][1],mult_result_i[47][0]}), .o_data(result_i[47*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000061_AdderTree0000000001(.i_data({mult_result_r[48][3],mult_result_r[48][2],mult_result_r[48][1],mult_result_r[48][0]}), .o_data(result_r[48*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000062_AdderTree0000000001(.i_data({mult_result_i[48][3],mult_result_i[48][2],mult_result_i[48][1],mult_result_i[48][0]}), .o_data(result_i[48*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000063_AdderTree0000000001(.i_data({mult_result_r[49][3],mult_result_r[49][2],mult_result_r[49][1],mult_result_r[49][0]}), .o_data(result_r[49*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000064_AdderTree0000000001(.i_data({mult_result_i[49][3],mult_result_i[49][2],mult_result_i[49][1],mult_result_i[49][0]}), .o_data(result_i[49*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000065_AdderTree0000000001(.i_data({mult_result_r[50][3],mult_result_r[50][2],mult_result_r[50][1],mult_result_r[50][0]}), .o_data(result_r[50*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000066_AdderTree0000000001(.i_data({mult_result_i[50][3],mult_result_i[50][2],mult_result_i[50][1],mult_result_i[50][0]}), .o_data(result_i[50*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000067_AdderTree0000000001(.i_data({mult_result_r[51][3],mult_result_r[51][2],mult_result_r[51][1],mult_result_r[51][0]}), .o_data(result_r[51*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000068_AdderTree0000000001(.i_data({mult_result_i[51][3],mult_result_i[51][2],mult_result_i[51][1],mult_result_i[51][0]}), .o_data(result_i[51*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000069_AdderTree0000000001(.i_data({mult_result_r[52][3],mult_result_r[52][2],mult_result_r[52][1],mult_result_r[52][0]}), .o_data(result_r[52*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000006A_AdderTree0000000001(.i_data({mult_result_i[52][3],mult_result_i[52][2],mult_result_i[52][1],mult_result_i[52][0]}), .o_data(result_i[52*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000006B_AdderTree0000000001(.i_data({mult_result_r[53][3],mult_result_r[53][2],mult_result_r[53][1],mult_result_r[53][0]}), .o_data(result_r[53*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000006C_AdderTree0000000001(.i_data({mult_result_i[53][3],mult_result_i[53][2],mult_result_i[53][1],mult_result_i[53][0]}), .o_data(result_i[53*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000006D_AdderTree0000000001(.i_data({mult_result_r[54][3],mult_result_r[54][2],mult_result_r[54][1],mult_result_r[54][0]}), .o_data(result_r[54*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000006E_AdderTree0000000001(.i_data({mult_result_i[54][3],mult_result_i[54][2],mult_result_i[54][1],mult_result_i[54][0]}), .o_data(result_i[54*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000006F_AdderTree0000000001(.i_data({mult_result_r[55][3],mult_result_r[55][2],mult_result_r[55][1],mult_result_r[55][0]}), .o_data(result_r[55*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000070_AdderTree0000000001(.i_data({mult_result_i[55][3],mult_result_i[55][2],mult_result_i[55][1],mult_result_i[55][0]}), .o_data(result_i[55*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000071_AdderTree0000000001(.i_data({mult_result_r[56][3],mult_result_r[56][2],mult_result_r[56][1],mult_result_r[56][0]}), .o_data(result_r[56*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000072_AdderTree0000000001(.i_data({mult_result_i[56][3],mult_result_i[56][2],mult_result_i[56][1],mult_result_i[56][0]}), .o_data(result_i[56*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000073_AdderTree0000000001(.i_data({mult_result_r[57][3],mult_result_r[57][2],mult_result_r[57][1],mult_result_r[57][0]}), .o_data(result_r[57*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000074_AdderTree0000000001(.i_data({mult_result_i[57][3],mult_result_i[57][2],mult_result_i[57][1],mult_result_i[57][0]}), .o_data(result_i[57*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000075_AdderTree0000000001(.i_data({mult_result_r[58][3],mult_result_r[58][2],mult_result_r[58][1],mult_result_r[58][0]}), .o_data(result_r[58*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000076_AdderTree0000000001(.i_data({mult_result_i[58][3],mult_result_i[58][2],mult_result_i[58][1],mult_result_i[58][0]}), .o_data(result_i[58*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000077_AdderTree0000000001(.i_data({mult_result_r[59][3],mult_result_r[59][2],mult_result_r[59][1],mult_result_r[59][0]}), .o_data(result_r[59*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000078_AdderTree0000000001(.i_data({mult_result_i[59][3],mult_result_i[59][2],mult_result_i[59][1],mult_result_i[59][0]}), .o_data(result_i[59*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000079_AdderTree0000000001(.i_data({mult_result_r[60][3],mult_result_r[60][2],mult_result_r[60][1],mult_result_r[60][0]}), .o_data(result_r[60*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000007A_AdderTree0000000001(.i_data({mult_result_i[60][3],mult_result_i[60][2],mult_result_i[60][1],mult_result_i[60][0]}), .o_data(result_i[60*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000007B_AdderTree0000000001(.i_data({mult_result_r[61][3],mult_result_r[61][2],mult_result_r[61][1],mult_result_r[61][0]}), .o_data(result_r[61*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000007C_AdderTree0000000001(.i_data({mult_result_i[61][3],mult_result_i[61][2],mult_result_i[61][1],mult_result_i[61][0]}), .o_data(result_i[61*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000007D_AdderTree0000000001(.i_data({mult_result_r[62][3],mult_result_r[62][2],mult_result_r[62][1],mult_result_r[62][0]}), .o_data(result_r[62*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000007E_AdderTree0000000001(.i_data({mult_result_i[62][3],mult_result_i[62][2],mult_result_i[62][1],mult_result_i[62][0]}), .o_data(result_i[62*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000007F_AdderTree0000000001(.i_data({mult_result_r[63][3],mult_result_r[63][2],mult_result_r[63][1],mult_result_r[63][0]}), .o_data(result_r[63*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000080_AdderTree0000000001(.i_data({mult_result_i[63][3],mult_result_i[63][2],mult_result_i[63][1],mult_result_i[63][0]}), .o_data(result_i[63*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000081_AdderTree0000000001(.i_data({mult_result_r[64][3],mult_result_r[64][2],mult_result_r[64][1],mult_result_r[64][0]}), .o_data(result_r[64*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000082_AdderTree0000000001(.i_data({mult_result_i[64][3],mult_result_i[64][2],mult_result_i[64][1],mult_result_i[64][0]}), .o_data(result_i[64*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000083_AdderTree0000000001(.i_data({mult_result_r[65][3],mult_result_r[65][2],mult_result_r[65][1],mult_result_r[65][0]}), .o_data(result_r[65*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000084_AdderTree0000000001(.i_data({mult_result_i[65][3],mult_result_i[65][2],mult_result_i[65][1],mult_result_i[65][0]}), .o_data(result_i[65*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000085_AdderTree0000000001(.i_data({mult_result_r[66][3],mult_result_r[66][2],mult_result_r[66][1],mult_result_r[66][0]}), .o_data(result_r[66*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000086_AdderTree0000000001(.i_data({mult_result_i[66][3],mult_result_i[66][2],mult_result_i[66][1],mult_result_i[66][0]}), .o_data(result_i[66*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000087_AdderTree0000000001(.i_data({mult_result_r[67][3],mult_result_r[67][2],mult_result_r[67][1],mult_result_r[67][0]}), .o_data(result_r[67*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000088_AdderTree0000000001(.i_data({mult_result_i[67][3],mult_result_i[67][2],mult_result_i[67][1],mult_result_i[67][0]}), .o_data(result_i[67*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000089_AdderTree0000000001(.i_data({mult_result_r[68][3],mult_result_r[68][2],mult_result_r[68][1],mult_result_r[68][0]}), .o_data(result_r[68*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000008A_AdderTree0000000001(.i_data({mult_result_i[68][3],mult_result_i[68][2],mult_result_i[68][1],mult_result_i[68][0]}), .o_data(result_i[68*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000008B_AdderTree0000000001(.i_data({mult_result_r[69][3],mult_result_r[69][2],mult_result_r[69][1],mult_result_r[69][0]}), .o_data(result_r[69*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000008C_AdderTree0000000001(.i_data({mult_result_i[69][3],mult_result_i[69][2],mult_result_i[69][1],mult_result_i[69][0]}), .o_data(result_i[69*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000008D_AdderTree0000000001(.i_data({mult_result_r[70][3],mult_result_r[70][2],mult_result_r[70][1],mult_result_r[70][0]}), .o_data(result_r[70*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000008E_AdderTree0000000001(.i_data({mult_result_i[70][3],mult_result_i[70][2],mult_result_i[70][1],mult_result_i[70][0]}), .o_data(result_i[70*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000008F_AdderTree0000000001(.i_data({mult_result_r[71][3],mult_result_r[71][2],mult_result_r[71][1],mult_result_r[71][0]}), .o_data(result_r[71*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000090_AdderTree0000000001(.i_data({mult_result_i[71][3],mult_result_i[71][2],mult_result_i[71][1],mult_result_i[71][0]}), .o_data(result_i[71*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000091_AdderTree0000000001(.i_data({mult_result_r[72][3],mult_result_r[72][2],mult_result_r[72][1],mult_result_r[72][0]}), .o_data(result_r[72*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000092_AdderTree0000000001(.i_data({mult_result_i[72][3],mult_result_i[72][2],mult_result_i[72][1],mult_result_i[72][0]}), .o_data(result_i[72*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000093_AdderTree0000000001(.i_data({mult_result_r[73][3],mult_result_r[73][2],mult_result_r[73][1],mult_result_r[73][0]}), .o_data(result_r[73*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000094_AdderTree0000000001(.i_data({mult_result_i[73][3],mult_result_i[73][2],mult_result_i[73][1],mult_result_i[73][0]}), .o_data(result_i[73*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000095_AdderTree0000000001(.i_data({mult_result_r[74][3],mult_result_r[74][2],mult_result_r[74][1],mult_result_r[74][0]}), .o_data(result_r[74*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000096_AdderTree0000000001(.i_data({mult_result_i[74][3],mult_result_i[74][2],mult_result_i[74][1],mult_result_i[74][0]}), .o_data(result_i[74*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000097_AdderTree0000000001(.i_data({mult_result_r[75][3],mult_result_r[75][2],mult_result_r[75][1],mult_result_r[75][0]}), .o_data(result_r[75*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000098_AdderTree0000000001(.i_data({mult_result_i[75][3],mult_result_i[75][2],mult_result_i[75][1],mult_result_i[75][0]}), .o_data(result_i[75*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000099_AdderTree0000000001(.i_data({mult_result_r[76][3],mult_result_r[76][2],mult_result_r[76][1],mult_result_r[76][0]}), .o_data(result_r[76*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000009A_AdderTree0000000001(.i_data({mult_result_i[76][3],mult_result_i[76][2],mult_result_i[76][1],mult_result_i[76][0]}), .o_data(result_i[76*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000009B_AdderTree0000000001(.i_data({mult_result_r[77][3],mult_result_r[77][2],mult_result_r[77][1],mult_result_r[77][0]}), .o_data(result_r[77*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000009C_AdderTree0000000001(.i_data({mult_result_i[77][3],mult_result_i[77][2],mult_result_i[77][1],mult_result_i[77][0]}), .o_data(result_i[77*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000009D_AdderTree0000000001(.i_data({mult_result_r[78][3],mult_result_r[78][2],mult_result_r[78][1],mult_result_r[78][0]}), .o_data(result_r[78*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000009E_AdderTree0000000001(.i_data({mult_result_i[78][3],mult_result_i[78][2],mult_result_i[78][1],mult_result_i[78][0]}), .o_data(result_i[78*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000009F_AdderTree0000000001(.i_data({mult_result_r[79][3],mult_result_r[79][2],mult_result_r[79][1],mult_result_r[79][0]}), .o_data(result_r[79*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000A0_AdderTree0000000001(.i_data({mult_result_i[79][3],mult_result_i[79][2],mult_result_i[79][1],mult_result_i[79][0]}), .o_data(result_i[79*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000A1_AdderTree0000000001(.i_data({mult_result_r[80][3],mult_result_r[80][2],mult_result_r[80][1],mult_result_r[80][0]}), .o_data(result_r[80*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000A2_AdderTree0000000001(.i_data({mult_result_i[80][3],mult_result_i[80][2],mult_result_i[80][1],mult_result_i[80][0]}), .o_data(result_i[80*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000A3_AdderTree0000000001(.i_data({mult_result_r[81][3],mult_result_r[81][2],mult_result_r[81][1],mult_result_r[81][0]}), .o_data(result_r[81*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000A4_AdderTree0000000001(.i_data({mult_result_i[81][3],mult_result_i[81][2],mult_result_i[81][1],mult_result_i[81][0]}), .o_data(result_i[81*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000A5_AdderTree0000000001(.i_data({mult_result_r[82][3],mult_result_r[82][2],mult_result_r[82][1],mult_result_r[82][0]}), .o_data(result_r[82*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000A6_AdderTree0000000001(.i_data({mult_result_i[82][3],mult_result_i[82][2],mult_result_i[82][1],mult_result_i[82][0]}), .o_data(result_i[82*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000A7_AdderTree0000000001(.i_data({mult_result_r[83][3],mult_result_r[83][2],mult_result_r[83][1],mult_result_r[83][0]}), .o_data(result_r[83*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000A8_AdderTree0000000001(.i_data({mult_result_i[83][3],mult_result_i[83][2],mult_result_i[83][1],mult_result_i[83][0]}), .o_data(result_i[83*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000A9_AdderTree0000000001(.i_data({mult_result_r[84][3],mult_result_r[84][2],mult_result_r[84][1],mult_result_r[84][0]}), .o_data(result_r[84*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000AA_AdderTree0000000001(.i_data({mult_result_i[84][3],mult_result_i[84][2],mult_result_i[84][1],mult_result_i[84][0]}), .o_data(result_i[84*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000AB_AdderTree0000000001(.i_data({mult_result_r[85][3],mult_result_r[85][2],mult_result_r[85][1],mult_result_r[85][0]}), .o_data(result_r[85*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000AC_AdderTree0000000001(.i_data({mult_result_i[85][3],mult_result_i[85][2],mult_result_i[85][1],mult_result_i[85][0]}), .o_data(result_i[85*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000AD_AdderTree0000000001(.i_data({mult_result_r[86][3],mult_result_r[86][2],mult_result_r[86][1],mult_result_r[86][0]}), .o_data(result_r[86*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000AE_AdderTree0000000001(.i_data({mult_result_i[86][3],mult_result_i[86][2],mult_result_i[86][1],mult_result_i[86][0]}), .o_data(result_i[86*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000AF_AdderTree0000000001(.i_data({mult_result_r[87][3],mult_result_r[87][2],mult_result_r[87][1],mult_result_r[87][0]}), .o_data(result_r[87*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000B0_AdderTree0000000001(.i_data({mult_result_i[87][3],mult_result_i[87][2],mult_result_i[87][1],mult_result_i[87][0]}), .o_data(result_i[87*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000B1_AdderTree0000000001(.i_data({mult_result_r[88][3],mult_result_r[88][2],mult_result_r[88][1],mult_result_r[88][0]}), .o_data(result_r[88*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000B2_AdderTree0000000001(.i_data({mult_result_i[88][3],mult_result_i[88][2],mult_result_i[88][1],mult_result_i[88][0]}), .o_data(result_i[88*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000B3_AdderTree0000000001(.i_data({mult_result_r[89][3],mult_result_r[89][2],mult_result_r[89][1],mult_result_r[89][0]}), .o_data(result_r[89*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000B4_AdderTree0000000001(.i_data({mult_result_i[89][3],mult_result_i[89][2],mult_result_i[89][1],mult_result_i[89][0]}), .o_data(result_i[89*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000B5_AdderTree0000000001(.i_data({mult_result_r[90][3],mult_result_r[90][2],mult_result_r[90][1],mult_result_r[90][0]}), .o_data(result_r[90*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000B6_AdderTree0000000001(.i_data({mult_result_i[90][3],mult_result_i[90][2],mult_result_i[90][1],mult_result_i[90][0]}), .o_data(result_i[90*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000B7_AdderTree0000000001(.i_data({mult_result_r[91][3],mult_result_r[91][2],mult_result_r[91][1],mult_result_r[91][0]}), .o_data(result_r[91*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000B8_AdderTree0000000001(.i_data({mult_result_i[91][3],mult_result_i[91][2],mult_result_i[91][1],mult_result_i[91][0]}), .o_data(result_i[91*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000B9_AdderTree0000000001(.i_data({mult_result_r[92][3],mult_result_r[92][2],mult_result_r[92][1],mult_result_r[92][0]}), .o_data(result_r[92*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000BA_AdderTree0000000001(.i_data({mult_result_i[92][3],mult_result_i[92][2],mult_result_i[92][1],mult_result_i[92][0]}), .o_data(result_i[92*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000BB_AdderTree0000000001(.i_data({mult_result_r[93][3],mult_result_r[93][2],mult_result_r[93][1],mult_result_r[93][0]}), .o_data(result_r[93*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000BC_AdderTree0000000001(.i_data({mult_result_i[93][3],mult_result_i[93][2],mult_result_i[93][1],mult_result_i[93][0]}), .o_data(result_i[93*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000BD_AdderTree0000000001(.i_data({mult_result_r[94][3],mult_result_r[94][2],mult_result_r[94][1],mult_result_r[94][0]}), .o_data(result_r[94*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000BE_AdderTree0000000001(.i_data({mult_result_i[94][3],mult_result_i[94][2],mult_result_i[94][1],mult_result_i[94][0]}), .o_data(result_i[94*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000BF_AdderTree0000000001(.i_data({mult_result_r[95][3],mult_result_r[95][2],mult_result_r[95][1],mult_result_r[95][0]}), .o_data(result_r[95*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000C0_AdderTree0000000001(.i_data({mult_result_i[95][3],mult_result_i[95][2],mult_result_i[95][1],mult_result_i[95][0]}), .o_data(result_i[95*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000C1_AdderTree0000000001(.i_data({mult_result_r[96][3],mult_result_r[96][2],mult_result_r[96][1],mult_result_r[96][0]}), .o_data(result_r[96*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000C2_AdderTree0000000001(.i_data({mult_result_i[96][3],mult_result_i[96][2],mult_result_i[96][1],mult_result_i[96][0]}), .o_data(result_i[96*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000C3_AdderTree0000000001(.i_data({mult_result_r[97][3],mult_result_r[97][2],mult_result_r[97][1],mult_result_r[97][0]}), .o_data(result_r[97*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000C4_AdderTree0000000001(.i_data({mult_result_i[97][3],mult_result_i[97][2],mult_result_i[97][1],mult_result_i[97][0]}), .o_data(result_i[97*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000C5_AdderTree0000000001(.i_data({mult_result_r[98][3],mult_result_r[98][2],mult_result_r[98][1],mult_result_r[98][0]}), .o_data(result_r[98*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000C6_AdderTree0000000001(.i_data({mult_result_i[98][3],mult_result_i[98][2],mult_result_i[98][1],mult_result_i[98][0]}), .o_data(result_i[98*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000C7_AdderTree0000000001(.i_data({mult_result_r[99][3],mult_result_r[99][2],mult_result_r[99][1],mult_result_r[99][0]}), .o_data(result_r[99*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000C8_AdderTree0000000001(.i_data({mult_result_i[99][3],mult_result_i[99][2],mult_result_i[99][1],mult_result_i[99][0]}), .o_data(result_i[99*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000C9_AdderTree0000000001(.i_data({mult_result_r[100][3],mult_result_r[100][2],mult_result_r[100][1],mult_result_r[100][0]}), .o_data(result_r[100*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000CA_AdderTree0000000001(.i_data({mult_result_i[100][3],mult_result_i[100][2],mult_result_i[100][1],mult_result_i[100][0]}), .o_data(result_i[100*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000CB_AdderTree0000000001(.i_data({mult_result_r[101][3],mult_result_r[101][2],mult_result_r[101][1],mult_result_r[101][0]}), .o_data(result_r[101*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000CC_AdderTree0000000001(.i_data({mult_result_i[101][3],mult_result_i[101][2],mult_result_i[101][1],mult_result_i[101][0]}), .o_data(result_i[101*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000CD_AdderTree0000000001(.i_data({mult_result_r[102][3],mult_result_r[102][2],mult_result_r[102][1],mult_result_r[102][0]}), .o_data(result_r[102*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000CE_AdderTree0000000001(.i_data({mult_result_i[102][3],mult_result_i[102][2],mult_result_i[102][1],mult_result_i[102][0]}), .o_data(result_i[102*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000CF_AdderTree0000000001(.i_data({mult_result_r[103][3],mult_result_r[103][2],mult_result_r[103][1],mult_result_r[103][0]}), .o_data(result_r[103*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000D0_AdderTree0000000001(.i_data({mult_result_i[103][3],mult_result_i[103][2],mult_result_i[103][1],mult_result_i[103][0]}), .o_data(result_i[103*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000D1_AdderTree0000000001(.i_data({mult_result_r[104][3],mult_result_r[104][2],mult_result_r[104][1],mult_result_r[104][0]}), .o_data(result_r[104*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000D2_AdderTree0000000001(.i_data({mult_result_i[104][3],mult_result_i[104][2],mult_result_i[104][1],mult_result_i[104][0]}), .o_data(result_i[104*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000D3_AdderTree0000000001(.i_data({mult_result_r[105][3],mult_result_r[105][2],mult_result_r[105][1],mult_result_r[105][0]}), .o_data(result_r[105*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000D4_AdderTree0000000001(.i_data({mult_result_i[105][3],mult_result_i[105][2],mult_result_i[105][1],mult_result_i[105][0]}), .o_data(result_i[105*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000D5_AdderTree0000000001(.i_data({mult_result_r[106][3],mult_result_r[106][2],mult_result_r[106][1],mult_result_r[106][0]}), .o_data(result_r[106*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000D6_AdderTree0000000001(.i_data({mult_result_i[106][3],mult_result_i[106][2],mult_result_i[106][1],mult_result_i[106][0]}), .o_data(result_i[106*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000D7_AdderTree0000000001(.i_data({mult_result_r[107][3],mult_result_r[107][2],mult_result_r[107][1],mult_result_r[107][0]}), .o_data(result_r[107*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000D8_AdderTree0000000001(.i_data({mult_result_i[107][3],mult_result_i[107][2],mult_result_i[107][1],mult_result_i[107][0]}), .o_data(result_i[107*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000D9_AdderTree0000000001(.i_data({mult_result_r[108][3],mult_result_r[108][2],mult_result_r[108][1],mult_result_r[108][0]}), .o_data(result_r[108*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000DA_AdderTree0000000001(.i_data({mult_result_i[108][3],mult_result_i[108][2],mult_result_i[108][1],mult_result_i[108][0]}), .o_data(result_i[108*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000DB_AdderTree0000000001(.i_data({mult_result_r[109][3],mult_result_r[109][2],mult_result_r[109][1],mult_result_r[109][0]}), .o_data(result_r[109*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000DC_AdderTree0000000001(.i_data({mult_result_i[109][3],mult_result_i[109][2],mult_result_i[109][1],mult_result_i[109][0]}), .o_data(result_i[109*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000DD_AdderTree0000000001(.i_data({mult_result_r[110][3],mult_result_r[110][2],mult_result_r[110][1],mult_result_r[110][0]}), .o_data(result_r[110*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000DE_AdderTree0000000001(.i_data({mult_result_i[110][3],mult_result_i[110][2],mult_result_i[110][1],mult_result_i[110][0]}), .o_data(result_i[110*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000DF_AdderTree0000000001(.i_data({mult_result_r[111][3],mult_result_r[111][2],mult_result_r[111][1],mult_result_r[111][0]}), .o_data(result_r[111*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000E0_AdderTree0000000001(.i_data({mult_result_i[111][3],mult_result_i[111][2],mult_result_i[111][1],mult_result_i[111][0]}), .o_data(result_i[111*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000E1_AdderTree0000000001(.i_data({mult_result_r[112][3],mult_result_r[112][2],mult_result_r[112][1],mult_result_r[112][0]}), .o_data(result_r[112*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000E2_AdderTree0000000001(.i_data({mult_result_i[112][3],mult_result_i[112][2],mult_result_i[112][1],mult_result_i[112][0]}), .o_data(result_i[112*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000E3_AdderTree0000000001(.i_data({mult_result_r[113][3],mult_result_r[113][2],mult_result_r[113][1],mult_result_r[113][0]}), .o_data(result_r[113*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000E4_AdderTree0000000001(.i_data({mult_result_i[113][3],mult_result_i[113][2],mult_result_i[113][1],mult_result_i[113][0]}), .o_data(result_i[113*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000E5_AdderTree0000000001(.i_data({mult_result_r[114][3],mult_result_r[114][2],mult_result_r[114][1],mult_result_r[114][0]}), .o_data(result_r[114*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000E6_AdderTree0000000001(.i_data({mult_result_i[114][3],mult_result_i[114][2],mult_result_i[114][1],mult_result_i[114][0]}), .o_data(result_i[114*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000E7_AdderTree0000000001(.i_data({mult_result_r[115][3],mult_result_r[115][2],mult_result_r[115][1],mult_result_r[115][0]}), .o_data(result_r[115*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000E8_AdderTree0000000001(.i_data({mult_result_i[115][3],mult_result_i[115][2],mult_result_i[115][1],mult_result_i[115][0]}), .o_data(result_i[115*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000E9_AdderTree0000000001(.i_data({mult_result_r[116][3],mult_result_r[116][2],mult_result_r[116][1],mult_result_r[116][0]}), .o_data(result_r[116*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000EA_AdderTree0000000001(.i_data({mult_result_i[116][3],mult_result_i[116][2],mult_result_i[116][1],mult_result_i[116][0]}), .o_data(result_i[116*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000EB_AdderTree0000000001(.i_data({mult_result_r[117][3],mult_result_r[117][2],mult_result_r[117][1],mult_result_r[117][0]}), .o_data(result_r[117*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000EC_AdderTree0000000001(.i_data({mult_result_i[117][3],mult_result_i[117][2],mult_result_i[117][1],mult_result_i[117][0]}), .o_data(result_i[117*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000ED_AdderTree0000000001(.i_data({mult_result_r[118][3],mult_result_r[118][2],mult_result_r[118][1],mult_result_r[118][0]}), .o_data(result_r[118*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000EE_AdderTree0000000001(.i_data({mult_result_i[118][3],mult_result_i[118][2],mult_result_i[118][1],mult_result_i[118][0]}), .o_data(result_i[118*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000EF_AdderTree0000000001(.i_data({mult_result_r[119][3],mult_result_r[119][2],mult_result_r[119][1],mult_result_r[119][0]}), .o_data(result_r[119*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000F0_AdderTree0000000001(.i_data({mult_result_i[119][3],mult_result_i[119][2],mult_result_i[119][1],mult_result_i[119][0]}), .o_data(result_i[119*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000F1_AdderTree0000000001(.i_data({mult_result_r[120][3],mult_result_r[120][2],mult_result_r[120][1],mult_result_r[120][0]}), .o_data(result_r[120*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000F2_AdderTree0000000001(.i_data({mult_result_i[120][3],mult_result_i[120][2],mult_result_i[120][1],mult_result_i[120][0]}), .o_data(result_i[120*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000F3_AdderTree0000000001(.i_data({mult_result_r[121][3],mult_result_r[121][2],mult_result_r[121][1],mult_result_r[121][0]}), .o_data(result_r[121*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000F4_AdderTree0000000001(.i_data({mult_result_i[121][3],mult_result_i[121][2],mult_result_i[121][1],mult_result_i[121][0]}), .o_data(result_i[121*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000F5_AdderTree0000000001(.i_data({mult_result_r[122][3],mult_result_r[122][2],mult_result_r[122][1],mult_result_r[122][0]}), .o_data(result_r[122*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000F6_AdderTree0000000001(.i_data({mult_result_i[122][3],mult_result_i[122][2],mult_result_i[122][1],mult_result_i[122][0]}), .o_data(result_i[122*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000F7_AdderTree0000000001(.i_data({mult_result_r[123][3],mult_result_r[123][2],mult_result_r[123][1],mult_result_r[123][0]}), .o_data(result_r[123*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000F8_AdderTree0000000001(.i_data({mult_result_i[123][3],mult_result_i[123][2],mult_result_i[123][1],mult_result_i[123][0]}), .o_data(result_i[123*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000F9_AdderTree0000000001(.i_data({mult_result_r[124][3],mult_result_r[124][2],mult_result_r[124][1],mult_result_r[124][0]}), .o_data(result_r[124*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000FA_AdderTree0000000001(.i_data({mult_result_i[124][3],mult_result_i[124][2],mult_result_i[124][1],mult_result_i[124][0]}), .o_data(result_i[124*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000FB_AdderTree0000000001(.i_data({mult_result_r[125][3],mult_result_r[125][2],mult_result_r[125][1],mult_result_r[125][0]}), .o_data(result_r[125*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000FC_AdderTree0000000001(.i_data({mult_result_i[125][3],mult_result_i[125][2],mult_result_i[125][1],mult_result_i[125][0]}), .o_data(result_i[125*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000FD_AdderTree0000000001(.i_data({mult_result_r[126][3],mult_result_r[126][2],mult_result_r[126][1],mult_result_r[126][0]}), .o_data(result_r[126*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000FE_AdderTree0000000001(.i_data({mult_result_i[126][3],mult_result_i[126][2],mult_result_i[126][1],mult_result_i[126][0]}), .o_data(result_i[126*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000000FF_AdderTree0000000001(.i_data({mult_result_r[127][3],mult_result_r[127][2],mult_result_r[127][1],mult_result_r[127][0]}), .o_data(result_r[127*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000100_AdderTree0000000001(.i_data({mult_result_i[127][3],mult_result_i[127][2],mult_result_i[127][1],mult_result_i[127][0]}), .o_data(result_i[127*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000101_AdderTree0000000001(.i_data({mult_result_r[128][3],mult_result_r[128][2],mult_result_r[128][1],mult_result_r[128][0]}), .o_data(result_r[128*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000102_AdderTree0000000001(.i_data({mult_result_i[128][3],mult_result_i[128][2],mult_result_i[128][1],mult_result_i[128][0]}), .o_data(result_i[128*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000103_AdderTree0000000001(.i_data({mult_result_r[129][3],mult_result_r[129][2],mult_result_r[129][1],mult_result_r[129][0]}), .o_data(result_r[129*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000104_AdderTree0000000001(.i_data({mult_result_i[129][3],mult_result_i[129][2],mult_result_i[129][1],mult_result_i[129][0]}), .o_data(result_i[129*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000105_AdderTree0000000001(.i_data({mult_result_r[130][3],mult_result_r[130][2],mult_result_r[130][1],mult_result_r[130][0]}), .o_data(result_r[130*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000106_AdderTree0000000001(.i_data({mult_result_i[130][3],mult_result_i[130][2],mult_result_i[130][1],mult_result_i[130][0]}), .o_data(result_i[130*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000107_AdderTree0000000001(.i_data({mult_result_r[131][3],mult_result_r[131][2],mult_result_r[131][1],mult_result_r[131][0]}), .o_data(result_r[131*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000108_AdderTree0000000001(.i_data({mult_result_i[131][3],mult_result_i[131][2],mult_result_i[131][1],mult_result_i[131][0]}), .o_data(result_i[131*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000109_AdderTree0000000001(.i_data({mult_result_r[132][3],mult_result_r[132][2],mult_result_r[132][1],mult_result_r[132][0]}), .o_data(result_r[132*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000010A_AdderTree0000000001(.i_data({mult_result_i[132][3],mult_result_i[132][2],mult_result_i[132][1],mult_result_i[132][0]}), .o_data(result_i[132*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000010B_AdderTree0000000001(.i_data({mult_result_r[133][3],mult_result_r[133][2],mult_result_r[133][1],mult_result_r[133][0]}), .o_data(result_r[133*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000010C_AdderTree0000000001(.i_data({mult_result_i[133][3],mult_result_i[133][2],mult_result_i[133][1],mult_result_i[133][0]}), .o_data(result_i[133*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000010D_AdderTree0000000001(.i_data({mult_result_r[134][3],mult_result_r[134][2],mult_result_r[134][1],mult_result_r[134][0]}), .o_data(result_r[134*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000010E_AdderTree0000000001(.i_data({mult_result_i[134][3],mult_result_i[134][2],mult_result_i[134][1],mult_result_i[134][0]}), .o_data(result_i[134*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000010F_AdderTree0000000001(.i_data({mult_result_r[135][3],mult_result_r[135][2],mult_result_r[135][1],mult_result_r[135][0]}), .o_data(result_r[135*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000110_AdderTree0000000001(.i_data({mult_result_i[135][3],mult_result_i[135][2],mult_result_i[135][1],mult_result_i[135][0]}), .o_data(result_i[135*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000111_AdderTree0000000001(.i_data({mult_result_r[136][3],mult_result_r[136][2],mult_result_r[136][1],mult_result_r[136][0]}), .o_data(result_r[136*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000112_AdderTree0000000001(.i_data({mult_result_i[136][3],mult_result_i[136][2],mult_result_i[136][1],mult_result_i[136][0]}), .o_data(result_i[136*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000113_AdderTree0000000001(.i_data({mult_result_r[137][3],mult_result_r[137][2],mult_result_r[137][1],mult_result_r[137][0]}), .o_data(result_r[137*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000114_AdderTree0000000001(.i_data({mult_result_i[137][3],mult_result_i[137][2],mult_result_i[137][1],mult_result_i[137][0]}), .o_data(result_i[137*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000115_AdderTree0000000001(.i_data({mult_result_r[138][3],mult_result_r[138][2],mult_result_r[138][1],mult_result_r[138][0]}), .o_data(result_r[138*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000116_AdderTree0000000001(.i_data({mult_result_i[138][3],mult_result_i[138][2],mult_result_i[138][1],mult_result_i[138][0]}), .o_data(result_i[138*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000117_AdderTree0000000001(.i_data({mult_result_r[139][3],mult_result_r[139][2],mult_result_r[139][1],mult_result_r[139][0]}), .o_data(result_r[139*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000118_AdderTree0000000001(.i_data({mult_result_i[139][3],mult_result_i[139][2],mult_result_i[139][1],mult_result_i[139][0]}), .o_data(result_i[139*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000119_AdderTree0000000001(.i_data({mult_result_r[140][3],mult_result_r[140][2],mult_result_r[140][1],mult_result_r[140][0]}), .o_data(result_r[140*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000011A_AdderTree0000000001(.i_data({mult_result_i[140][3],mult_result_i[140][2],mult_result_i[140][1],mult_result_i[140][0]}), .o_data(result_i[140*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000011B_AdderTree0000000001(.i_data({mult_result_r[141][3],mult_result_r[141][2],mult_result_r[141][1],mult_result_r[141][0]}), .o_data(result_r[141*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000011C_AdderTree0000000001(.i_data({mult_result_i[141][3],mult_result_i[141][2],mult_result_i[141][1],mult_result_i[141][0]}), .o_data(result_i[141*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000011D_AdderTree0000000001(.i_data({mult_result_r[142][3],mult_result_r[142][2],mult_result_r[142][1],mult_result_r[142][0]}), .o_data(result_r[142*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000011E_AdderTree0000000001(.i_data({mult_result_i[142][3],mult_result_i[142][2],mult_result_i[142][1],mult_result_i[142][0]}), .o_data(result_i[142*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000011F_AdderTree0000000001(.i_data({mult_result_r[143][3],mult_result_r[143][2],mult_result_r[143][1],mult_result_r[143][0]}), .o_data(result_r[143*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000120_AdderTree0000000001(.i_data({mult_result_i[143][3],mult_result_i[143][2],mult_result_i[143][1],mult_result_i[143][0]}), .o_data(result_i[143*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000121_AdderTree0000000001(.i_data({mult_result_r[144][3],mult_result_r[144][2],mult_result_r[144][1],mult_result_r[144][0]}), .o_data(result_r[144*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000122_AdderTree0000000001(.i_data({mult_result_i[144][3],mult_result_i[144][2],mult_result_i[144][1],mult_result_i[144][0]}), .o_data(result_i[144*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000123_AdderTree0000000001(.i_data({mult_result_r[145][3],mult_result_r[145][2],mult_result_r[145][1],mult_result_r[145][0]}), .o_data(result_r[145*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000124_AdderTree0000000001(.i_data({mult_result_i[145][3],mult_result_i[145][2],mult_result_i[145][1],mult_result_i[145][0]}), .o_data(result_i[145*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000125_AdderTree0000000001(.i_data({mult_result_r[146][3],mult_result_r[146][2],mult_result_r[146][1],mult_result_r[146][0]}), .o_data(result_r[146*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000126_AdderTree0000000001(.i_data({mult_result_i[146][3],mult_result_i[146][2],mult_result_i[146][1],mult_result_i[146][0]}), .o_data(result_i[146*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000127_AdderTree0000000001(.i_data({mult_result_r[147][3],mult_result_r[147][2],mult_result_r[147][1],mult_result_r[147][0]}), .o_data(result_r[147*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000128_AdderTree0000000001(.i_data({mult_result_i[147][3],mult_result_i[147][2],mult_result_i[147][1],mult_result_i[147][0]}), .o_data(result_i[147*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000129_AdderTree0000000001(.i_data({mult_result_r[148][3],mult_result_r[148][2],mult_result_r[148][1],mult_result_r[148][0]}), .o_data(result_r[148*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000012A_AdderTree0000000001(.i_data({mult_result_i[148][3],mult_result_i[148][2],mult_result_i[148][1],mult_result_i[148][0]}), .o_data(result_i[148*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000012B_AdderTree0000000001(.i_data({mult_result_r[149][3],mult_result_r[149][2],mult_result_r[149][1],mult_result_r[149][0]}), .o_data(result_r[149*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000012C_AdderTree0000000001(.i_data({mult_result_i[149][3],mult_result_i[149][2],mult_result_i[149][1],mult_result_i[149][0]}), .o_data(result_i[149*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000012D_AdderTree0000000001(.i_data({mult_result_r[150][3],mult_result_r[150][2],mult_result_r[150][1],mult_result_r[150][0]}), .o_data(result_r[150*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000012E_AdderTree0000000001(.i_data({mult_result_i[150][3],mult_result_i[150][2],mult_result_i[150][1],mult_result_i[150][0]}), .o_data(result_i[150*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000012F_AdderTree0000000001(.i_data({mult_result_r[151][3],mult_result_r[151][2],mult_result_r[151][1],mult_result_r[151][0]}), .o_data(result_r[151*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000130_AdderTree0000000001(.i_data({mult_result_i[151][3],mult_result_i[151][2],mult_result_i[151][1],mult_result_i[151][0]}), .o_data(result_i[151*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000131_AdderTree0000000001(.i_data({mult_result_r[152][3],mult_result_r[152][2],mult_result_r[152][1],mult_result_r[152][0]}), .o_data(result_r[152*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000132_AdderTree0000000001(.i_data({mult_result_i[152][3],mult_result_i[152][2],mult_result_i[152][1],mult_result_i[152][0]}), .o_data(result_i[152*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000133_AdderTree0000000001(.i_data({mult_result_r[153][3],mult_result_r[153][2],mult_result_r[153][1],mult_result_r[153][0]}), .o_data(result_r[153*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000134_AdderTree0000000001(.i_data({mult_result_i[153][3],mult_result_i[153][2],mult_result_i[153][1],mult_result_i[153][0]}), .o_data(result_i[153*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000135_AdderTree0000000001(.i_data({mult_result_r[154][3],mult_result_r[154][2],mult_result_r[154][1],mult_result_r[154][0]}), .o_data(result_r[154*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000136_AdderTree0000000001(.i_data({mult_result_i[154][3],mult_result_i[154][2],mult_result_i[154][1],mult_result_i[154][0]}), .o_data(result_i[154*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000137_AdderTree0000000001(.i_data({mult_result_r[155][3],mult_result_r[155][2],mult_result_r[155][1],mult_result_r[155][0]}), .o_data(result_r[155*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000138_AdderTree0000000001(.i_data({mult_result_i[155][3],mult_result_i[155][2],mult_result_i[155][1],mult_result_i[155][0]}), .o_data(result_i[155*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000139_AdderTree0000000001(.i_data({mult_result_r[156][3],mult_result_r[156][2],mult_result_r[156][1],mult_result_r[156][0]}), .o_data(result_r[156*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000013A_AdderTree0000000001(.i_data({mult_result_i[156][3],mult_result_i[156][2],mult_result_i[156][1],mult_result_i[156][0]}), .o_data(result_i[156*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000013B_AdderTree0000000001(.i_data({mult_result_r[157][3],mult_result_r[157][2],mult_result_r[157][1],mult_result_r[157][0]}), .o_data(result_r[157*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000013C_AdderTree0000000001(.i_data({mult_result_i[157][3],mult_result_i[157][2],mult_result_i[157][1],mult_result_i[157][0]}), .o_data(result_i[157*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000013D_AdderTree0000000001(.i_data({mult_result_r[158][3],mult_result_r[158][2],mult_result_r[158][1],mult_result_r[158][0]}), .o_data(result_r[158*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000013E_AdderTree0000000001(.i_data({mult_result_i[158][3],mult_result_i[158][2],mult_result_i[158][1],mult_result_i[158][0]}), .o_data(result_i[158*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000013F_AdderTree0000000001(.i_data({mult_result_r[159][3],mult_result_r[159][2],mult_result_r[159][1],mult_result_r[159][0]}), .o_data(result_r[159*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000140_AdderTree0000000001(.i_data({mult_result_i[159][3],mult_result_i[159][2],mult_result_i[159][1],mult_result_i[159][0]}), .o_data(result_i[159*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000141_AdderTree0000000001(.i_data({mult_result_r[160][3],mult_result_r[160][2],mult_result_r[160][1],mult_result_r[160][0]}), .o_data(result_r[160*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000142_AdderTree0000000001(.i_data({mult_result_i[160][3],mult_result_i[160][2],mult_result_i[160][1],mult_result_i[160][0]}), .o_data(result_i[160*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000143_AdderTree0000000001(.i_data({mult_result_r[161][3],mult_result_r[161][2],mult_result_r[161][1],mult_result_r[161][0]}), .o_data(result_r[161*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000144_AdderTree0000000001(.i_data({mult_result_i[161][3],mult_result_i[161][2],mult_result_i[161][1],mult_result_i[161][0]}), .o_data(result_i[161*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000145_AdderTree0000000001(.i_data({mult_result_r[162][3],mult_result_r[162][2],mult_result_r[162][1],mult_result_r[162][0]}), .o_data(result_r[162*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000146_AdderTree0000000001(.i_data({mult_result_i[162][3],mult_result_i[162][2],mult_result_i[162][1],mult_result_i[162][0]}), .o_data(result_i[162*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000147_AdderTree0000000001(.i_data({mult_result_r[163][3],mult_result_r[163][2],mult_result_r[163][1],mult_result_r[163][0]}), .o_data(result_r[163*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000148_AdderTree0000000001(.i_data({mult_result_i[163][3],mult_result_i[163][2],mult_result_i[163][1],mult_result_i[163][0]}), .o_data(result_i[163*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000149_AdderTree0000000001(.i_data({mult_result_r[164][3],mult_result_r[164][2],mult_result_r[164][1],mult_result_r[164][0]}), .o_data(result_r[164*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000014A_AdderTree0000000001(.i_data({mult_result_i[164][3],mult_result_i[164][2],mult_result_i[164][1],mult_result_i[164][0]}), .o_data(result_i[164*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000014B_AdderTree0000000001(.i_data({mult_result_r[165][3],mult_result_r[165][2],mult_result_r[165][1],mult_result_r[165][0]}), .o_data(result_r[165*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000014C_AdderTree0000000001(.i_data({mult_result_i[165][3],mult_result_i[165][2],mult_result_i[165][1],mult_result_i[165][0]}), .o_data(result_i[165*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000014D_AdderTree0000000001(.i_data({mult_result_r[166][3],mult_result_r[166][2],mult_result_r[166][1],mult_result_r[166][0]}), .o_data(result_r[166*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000014E_AdderTree0000000001(.i_data({mult_result_i[166][3],mult_result_i[166][2],mult_result_i[166][1],mult_result_i[166][0]}), .o_data(result_i[166*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000014F_AdderTree0000000001(.i_data({mult_result_r[167][3],mult_result_r[167][2],mult_result_r[167][1],mult_result_r[167][0]}), .o_data(result_r[167*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000150_AdderTree0000000001(.i_data({mult_result_i[167][3],mult_result_i[167][2],mult_result_i[167][1],mult_result_i[167][0]}), .o_data(result_i[167*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000151_AdderTree0000000001(.i_data({mult_result_r[168][3],mult_result_r[168][2],mult_result_r[168][1],mult_result_r[168][0]}), .o_data(result_r[168*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000152_AdderTree0000000001(.i_data({mult_result_i[168][3],mult_result_i[168][2],mult_result_i[168][1],mult_result_i[168][0]}), .o_data(result_i[168*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000153_AdderTree0000000001(.i_data({mult_result_r[169][3],mult_result_r[169][2],mult_result_r[169][1],mult_result_r[169][0]}), .o_data(result_r[169*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000154_AdderTree0000000001(.i_data({mult_result_i[169][3],mult_result_i[169][2],mult_result_i[169][1],mult_result_i[169][0]}), .o_data(result_i[169*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000155_AdderTree0000000001(.i_data({mult_result_r[170][3],mult_result_r[170][2],mult_result_r[170][1],mult_result_r[170][0]}), .o_data(result_r[170*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000156_AdderTree0000000001(.i_data({mult_result_i[170][3],mult_result_i[170][2],mult_result_i[170][1],mult_result_i[170][0]}), .o_data(result_i[170*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000157_AdderTree0000000001(.i_data({mult_result_r[171][3],mult_result_r[171][2],mult_result_r[171][1],mult_result_r[171][0]}), .o_data(result_r[171*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000158_AdderTree0000000001(.i_data({mult_result_i[171][3],mult_result_i[171][2],mult_result_i[171][1],mult_result_i[171][0]}), .o_data(result_i[171*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000159_AdderTree0000000001(.i_data({mult_result_r[172][3],mult_result_r[172][2],mult_result_r[172][1],mult_result_r[172][0]}), .o_data(result_r[172*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000015A_AdderTree0000000001(.i_data({mult_result_i[172][3],mult_result_i[172][2],mult_result_i[172][1],mult_result_i[172][0]}), .o_data(result_i[172*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000015B_AdderTree0000000001(.i_data({mult_result_r[173][3],mult_result_r[173][2],mult_result_r[173][1],mult_result_r[173][0]}), .o_data(result_r[173*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000015C_AdderTree0000000001(.i_data({mult_result_i[173][3],mult_result_i[173][2],mult_result_i[173][1],mult_result_i[173][0]}), .o_data(result_i[173*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000015D_AdderTree0000000001(.i_data({mult_result_r[174][3],mult_result_r[174][2],mult_result_r[174][1],mult_result_r[174][0]}), .o_data(result_r[174*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000015E_AdderTree0000000001(.i_data({mult_result_i[174][3],mult_result_i[174][2],mult_result_i[174][1],mult_result_i[174][0]}), .o_data(result_i[174*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000015F_AdderTree0000000001(.i_data({mult_result_r[175][3],mult_result_r[175][2],mult_result_r[175][1],mult_result_r[175][0]}), .o_data(result_r[175*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000160_AdderTree0000000001(.i_data({mult_result_i[175][3],mult_result_i[175][2],mult_result_i[175][1],mult_result_i[175][0]}), .o_data(result_i[175*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000161_AdderTree0000000001(.i_data({mult_result_r[176][3],mult_result_r[176][2],mult_result_r[176][1],mult_result_r[176][0]}), .o_data(result_r[176*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000162_AdderTree0000000001(.i_data({mult_result_i[176][3],mult_result_i[176][2],mult_result_i[176][1],mult_result_i[176][0]}), .o_data(result_i[176*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000163_AdderTree0000000001(.i_data({mult_result_r[177][3],mult_result_r[177][2],mult_result_r[177][1],mult_result_r[177][0]}), .o_data(result_r[177*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000164_AdderTree0000000001(.i_data({mult_result_i[177][3],mult_result_i[177][2],mult_result_i[177][1],mult_result_i[177][0]}), .o_data(result_i[177*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000165_AdderTree0000000001(.i_data({mult_result_r[178][3],mult_result_r[178][2],mult_result_r[178][1],mult_result_r[178][0]}), .o_data(result_r[178*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000166_AdderTree0000000001(.i_data({mult_result_i[178][3],mult_result_i[178][2],mult_result_i[178][1],mult_result_i[178][0]}), .o_data(result_i[178*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000167_AdderTree0000000001(.i_data({mult_result_r[179][3],mult_result_r[179][2],mult_result_r[179][1],mult_result_r[179][0]}), .o_data(result_r[179*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000168_AdderTree0000000001(.i_data({mult_result_i[179][3],mult_result_i[179][2],mult_result_i[179][1],mult_result_i[179][0]}), .o_data(result_i[179*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000169_AdderTree0000000001(.i_data({mult_result_r[180][3],mult_result_r[180][2],mult_result_r[180][1],mult_result_r[180][0]}), .o_data(result_r[180*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000016A_AdderTree0000000001(.i_data({mult_result_i[180][3],mult_result_i[180][2],mult_result_i[180][1],mult_result_i[180][0]}), .o_data(result_i[180*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000016B_AdderTree0000000001(.i_data({mult_result_r[181][3],mult_result_r[181][2],mult_result_r[181][1],mult_result_r[181][0]}), .o_data(result_r[181*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000016C_AdderTree0000000001(.i_data({mult_result_i[181][3],mult_result_i[181][2],mult_result_i[181][1],mult_result_i[181][0]}), .o_data(result_i[181*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000016D_AdderTree0000000001(.i_data({mult_result_r[182][3],mult_result_r[182][2],mult_result_r[182][1],mult_result_r[182][0]}), .o_data(result_r[182*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000016E_AdderTree0000000001(.i_data({mult_result_i[182][3],mult_result_i[182][2],mult_result_i[182][1],mult_result_i[182][0]}), .o_data(result_i[182*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000016F_AdderTree0000000001(.i_data({mult_result_r[183][3],mult_result_r[183][2],mult_result_r[183][1],mult_result_r[183][0]}), .o_data(result_r[183*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000170_AdderTree0000000001(.i_data({mult_result_i[183][3],mult_result_i[183][2],mult_result_i[183][1],mult_result_i[183][0]}), .o_data(result_i[183*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000171_AdderTree0000000001(.i_data({mult_result_r[184][3],mult_result_r[184][2],mult_result_r[184][1],mult_result_r[184][0]}), .o_data(result_r[184*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000172_AdderTree0000000001(.i_data({mult_result_i[184][3],mult_result_i[184][2],mult_result_i[184][1],mult_result_i[184][0]}), .o_data(result_i[184*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000173_AdderTree0000000001(.i_data({mult_result_r[185][3],mult_result_r[185][2],mult_result_r[185][1],mult_result_r[185][0]}), .o_data(result_r[185*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000174_AdderTree0000000001(.i_data({mult_result_i[185][3],mult_result_i[185][2],mult_result_i[185][1],mult_result_i[185][0]}), .o_data(result_i[185*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000175_AdderTree0000000001(.i_data({mult_result_r[186][3],mult_result_r[186][2],mult_result_r[186][1],mult_result_r[186][0]}), .o_data(result_r[186*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000176_AdderTree0000000001(.i_data({mult_result_i[186][3],mult_result_i[186][2],mult_result_i[186][1],mult_result_i[186][0]}), .o_data(result_i[186*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000177_AdderTree0000000001(.i_data({mult_result_r[187][3],mult_result_r[187][2],mult_result_r[187][1],mult_result_r[187][0]}), .o_data(result_r[187*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000178_AdderTree0000000001(.i_data({mult_result_i[187][3],mult_result_i[187][2],mult_result_i[187][1],mult_result_i[187][0]}), .o_data(result_i[187*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000179_AdderTree0000000001(.i_data({mult_result_r[188][3],mult_result_r[188][2],mult_result_r[188][1],mult_result_r[188][0]}), .o_data(result_r[188*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000017A_AdderTree0000000001(.i_data({mult_result_i[188][3],mult_result_i[188][2],mult_result_i[188][1],mult_result_i[188][0]}), .o_data(result_i[188*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000017B_AdderTree0000000001(.i_data({mult_result_r[189][3],mult_result_r[189][2],mult_result_r[189][1],mult_result_r[189][0]}), .o_data(result_r[189*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000017C_AdderTree0000000001(.i_data({mult_result_i[189][3],mult_result_i[189][2],mult_result_i[189][1],mult_result_i[189][0]}), .o_data(result_i[189*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000017D_AdderTree0000000001(.i_data({mult_result_r[190][3],mult_result_r[190][2],mult_result_r[190][1],mult_result_r[190][0]}), .o_data(result_r[190*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000017E_AdderTree0000000001(.i_data({mult_result_i[190][3],mult_result_i[190][2],mult_result_i[190][1],mult_result_i[190][0]}), .o_data(result_i[190*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000017F_AdderTree0000000001(.i_data({mult_result_r[191][3],mult_result_r[191][2],mult_result_r[191][1],mult_result_r[191][0]}), .o_data(result_r[191*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000180_AdderTree0000000001(.i_data({mult_result_i[191][3],mult_result_i[191][2],mult_result_i[191][1],mult_result_i[191][0]}), .o_data(result_i[191*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000181_AdderTree0000000001(.i_data({mult_result_r[192][3],mult_result_r[192][2],mult_result_r[192][1],mult_result_r[192][0]}), .o_data(result_r[192*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000182_AdderTree0000000001(.i_data({mult_result_i[192][3],mult_result_i[192][2],mult_result_i[192][1],mult_result_i[192][0]}), .o_data(result_i[192*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000183_AdderTree0000000001(.i_data({mult_result_r[193][3],mult_result_r[193][2],mult_result_r[193][1],mult_result_r[193][0]}), .o_data(result_r[193*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000184_AdderTree0000000001(.i_data({mult_result_i[193][3],mult_result_i[193][2],mult_result_i[193][1],mult_result_i[193][0]}), .o_data(result_i[193*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000185_AdderTree0000000001(.i_data({mult_result_r[194][3],mult_result_r[194][2],mult_result_r[194][1],mult_result_r[194][0]}), .o_data(result_r[194*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000186_AdderTree0000000001(.i_data({mult_result_i[194][3],mult_result_i[194][2],mult_result_i[194][1],mult_result_i[194][0]}), .o_data(result_i[194*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000187_AdderTree0000000001(.i_data({mult_result_r[195][3],mult_result_r[195][2],mult_result_r[195][1],mult_result_r[195][0]}), .o_data(result_r[195*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000188_AdderTree0000000001(.i_data({mult_result_i[195][3],mult_result_i[195][2],mult_result_i[195][1],mult_result_i[195][0]}), .o_data(result_i[195*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000189_AdderTree0000000001(.i_data({mult_result_r[196][3],mult_result_r[196][2],mult_result_r[196][1],mult_result_r[196][0]}), .o_data(result_r[196*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000018A_AdderTree0000000001(.i_data({mult_result_i[196][3],mult_result_i[196][2],mult_result_i[196][1],mult_result_i[196][0]}), .o_data(result_i[196*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000018B_AdderTree0000000001(.i_data({mult_result_r[197][3],mult_result_r[197][2],mult_result_r[197][1],mult_result_r[197][0]}), .o_data(result_r[197*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000018C_AdderTree0000000001(.i_data({mult_result_i[197][3],mult_result_i[197][2],mult_result_i[197][1],mult_result_i[197][0]}), .o_data(result_i[197*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000018D_AdderTree0000000001(.i_data({mult_result_r[198][3],mult_result_r[198][2],mult_result_r[198][1],mult_result_r[198][0]}), .o_data(result_r[198*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000018E_AdderTree0000000001(.i_data({mult_result_i[198][3],mult_result_i[198][2],mult_result_i[198][1],mult_result_i[198][0]}), .o_data(result_i[198*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000018F_AdderTree0000000001(.i_data({mult_result_r[199][3],mult_result_r[199][2],mult_result_r[199][1],mult_result_r[199][0]}), .o_data(result_r[199*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000190_AdderTree0000000001(.i_data({mult_result_i[199][3],mult_result_i[199][2],mult_result_i[199][1],mult_result_i[199][0]}), .o_data(result_i[199*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000191_AdderTree0000000001(.i_data({mult_result_r[200][3],mult_result_r[200][2],mult_result_r[200][1],mult_result_r[200][0]}), .o_data(result_r[200*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000192_AdderTree0000000001(.i_data({mult_result_i[200][3],mult_result_i[200][2],mult_result_i[200][1],mult_result_i[200][0]}), .o_data(result_i[200*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000193_AdderTree0000000001(.i_data({mult_result_r[201][3],mult_result_r[201][2],mult_result_r[201][1],mult_result_r[201][0]}), .o_data(result_r[201*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000194_AdderTree0000000001(.i_data({mult_result_i[201][3],mult_result_i[201][2],mult_result_i[201][1],mult_result_i[201][0]}), .o_data(result_i[201*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000195_AdderTree0000000001(.i_data({mult_result_r[202][3],mult_result_r[202][2],mult_result_r[202][1],mult_result_r[202][0]}), .o_data(result_r[202*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000196_AdderTree0000000001(.i_data({mult_result_i[202][3],mult_result_i[202][2],mult_result_i[202][1],mult_result_i[202][0]}), .o_data(result_i[202*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000197_AdderTree0000000001(.i_data({mult_result_r[203][3],mult_result_r[203][2],mult_result_r[203][1],mult_result_r[203][0]}), .o_data(result_r[203*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000198_AdderTree0000000001(.i_data({mult_result_i[203][3],mult_result_i[203][2],mult_result_i[203][1],mult_result_i[203][0]}), .o_data(result_i[203*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000199_AdderTree0000000001(.i_data({mult_result_r[204][3],mult_result_r[204][2],mult_result_r[204][1],mult_result_r[204][0]}), .o_data(result_r[204*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000019A_AdderTree0000000001(.i_data({mult_result_i[204][3],mult_result_i[204][2],mult_result_i[204][1],mult_result_i[204][0]}), .o_data(result_i[204*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000019B_AdderTree0000000001(.i_data({mult_result_r[205][3],mult_result_r[205][2],mult_result_r[205][1],mult_result_r[205][0]}), .o_data(result_r[205*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000019C_AdderTree0000000001(.i_data({mult_result_i[205][3],mult_result_i[205][2],mult_result_i[205][1],mult_result_i[205][0]}), .o_data(result_i[205*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000019D_AdderTree0000000001(.i_data({mult_result_r[206][3],mult_result_r[206][2],mult_result_r[206][1],mult_result_r[206][0]}), .o_data(result_r[206*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000019E_AdderTree0000000001(.i_data({mult_result_i[206][3],mult_result_i[206][2],mult_result_i[206][1],mult_result_i[206][0]}), .o_data(result_i[206*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_000000019F_AdderTree0000000001(.i_data({mult_result_r[207][3],mult_result_r[207][2],mult_result_r[207][1],mult_result_r[207][0]}), .o_data(result_r[207*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001A0_AdderTree0000000001(.i_data({mult_result_i[207][3],mult_result_i[207][2],mult_result_i[207][1],mult_result_i[207][0]}), .o_data(result_i[207*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001A1_AdderTree0000000001(.i_data({mult_result_r[208][3],mult_result_r[208][2],mult_result_r[208][1],mult_result_r[208][0]}), .o_data(result_r[208*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001A2_AdderTree0000000001(.i_data({mult_result_i[208][3],mult_result_i[208][2],mult_result_i[208][1],mult_result_i[208][0]}), .o_data(result_i[208*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001A3_AdderTree0000000001(.i_data({mult_result_r[209][3],mult_result_r[209][2],mult_result_r[209][1],mult_result_r[209][0]}), .o_data(result_r[209*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001A4_AdderTree0000000001(.i_data({mult_result_i[209][3],mult_result_i[209][2],mult_result_i[209][1],mult_result_i[209][0]}), .o_data(result_i[209*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001A5_AdderTree0000000001(.i_data({mult_result_r[210][3],mult_result_r[210][2],mult_result_r[210][1],mult_result_r[210][0]}), .o_data(result_r[210*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001A6_AdderTree0000000001(.i_data({mult_result_i[210][3],mult_result_i[210][2],mult_result_i[210][1],mult_result_i[210][0]}), .o_data(result_i[210*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001A7_AdderTree0000000001(.i_data({mult_result_r[211][3],mult_result_r[211][2],mult_result_r[211][1],mult_result_r[211][0]}), .o_data(result_r[211*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001A8_AdderTree0000000001(.i_data({mult_result_i[211][3],mult_result_i[211][2],mult_result_i[211][1],mult_result_i[211][0]}), .o_data(result_i[211*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001A9_AdderTree0000000001(.i_data({mult_result_r[212][3],mult_result_r[212][2],mult_result_r[212][1],mult_result_r[212][0]}), .o_data(result_r[212*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001AA_AdderTree0000000001(.i_data({mult_result_i[212][3],mult_result_i[212][2],mult_result_i[212][1],mult_result_i[212][0]}), .o_data(result_i[212*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001AB_AdderTree0000000001(.i_data({mult_result_r[213][3],mult_result_r[213][2],mult_result_r[213][1],mult_result_r[213][0]}), .o_data(result_r[213*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001AC_AdderTree0000000001(.i_data({mult_result_i[213][3],mult_result_i[213][2],mult_result_i[213][1],mult_result_i[213][0]}), .o_data(result_i[213*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001AD_AdderTree0000000001(.i_data({mult_result_r[214][3],mult_result_r[214][2],mult_result_r[214][1],mult_result_r[214][0]}), .o_data(result_r[214*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001AE_AdderTree0000000001(.i_data({mult_result_i[214][3],mult_result_i[214][2],mult_result_i[214][1],mult_result_i[214][0]}), .o_data(result_i[214*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001AF_AdderTree0000000001(.i_data({mult_result_r[215][3],mult_result_r[215][2],mult_result_r[215][1],mult_result_r[215][0]}), .o_data(result_r[215*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001B0_AdderTree0000000001(.i_data({mult_result_i[215][3],mult_result_i[215][2],mult_result_i[215][1],mult_result_i[215][0]}), .o_data(result_i[215*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001B1_AdderTree0000000001(.i_data({mult_result_r[216][3],mult_result_r[216][2],mult_result_r[216][1],mult_result_r[216][0]}), .o_data(result_r[216*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001B2_AdderTree0000000001(.i_data({mult_result_i[216][3],mult_result_i[216][2],mult_result_i[216][1],mult_result_i[216][0]}), .o_data(result_i[216*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001B3_AdderTree0000000001(.i_data({mult_result_r[217][3],mult_result_r[217][2],mult_result_r[217][1],mult_result_r[217][0]}), .o_data(result_r[217*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001B4_AdderTree0000000001(.i_data({mult_result_i[217][3],mult_result_i[217][2],mult_result_i[217][1],mult_result_i[217][0]}), .o_data(result_i[217*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001B5_AdderTree0000000001(.i_data({mult_result_r[218][3],mult_result_r[218][2],mult_result_r[218][1],mult_result_r[218][0]}), .o_data(result_r[218*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001B6_AdderTree0000000001(.i_data({mult_result_i[218][3],mult_result_i[218][2],mult_result_i[218][1],mult_result_i[218][0]}), .o_data(result_i[218*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001B7_AdderTree0000000001(.i_data({mult_result_r[219][3],mult_result_r[219][2],mult_result_r[219][1],mult_result_r[219][0]}), .o_data(result_r[219*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001B8_AdderTree0000000001(.i_data({mult_result_i[219][3],mult_result_i[219][2],mult_result_i[219][1],mult_result_i[219][0]}), .o_data(result_i[219*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001B9_AdderTree0000000001(.i_data({mult_result_r[220][3],mult_result_r[220][2],mult_result_r[220][1],mult_result_r[220][0]}), .o_data(result_r[220*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001BA_AdderTree0000000001(.i_data({mult_result_i[220][3],mult_result_i[220][2],mult_result_i[220][1],mult_result_i[220][0]}), .o_data(result_i[220*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001BB_AdderTree0000000001(.i_data({mult_result_r[221][3],mult_result_r[221][2],mult_result_r[221][1],mult_result_r[221][0]}), .o_data(result_r[221*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001BC_AdderTree0000000001(.i_data({mult_result_i[221][3],mult_result_i[221][2],mult_result_i[221][1],mult_result_i[221][0]}), .o_data(result_i[221*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001BD_AdderTree0000000001(.i_data({mult_result_r[222][3],mult_result_r[222][2],mult_result_r[222][1],mult_result_r[222][0]}), .o_data(result_r[222*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001BE_AdderTree0000000001(.i_data({mult_result_i[222][3],mult_result_i[222][2],mult_result_i[222][1],mult_result_i[222][0]}), .o_data(result_i[222*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001BF_AdderTree0000000001(.i_data({mult_result_r[223][3],mult_result_r[223][2],mult_result_r[223][1],mult_result_r[223][0]}), .o_data(result_r[223*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001C0_AdderTree0000000001(.i_data({mult_result_i[223][3],mult_result_i[223][2],mult_result_i[223][1],mult_result_i[223][0]}), .o_data(result_i[223*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001C1_AdderTree0000000001(.i_data({mult_result_r[224][3],mult_result_r[224][2],mult_result_r[224][1],mult_result_r[224][0]}), .o_data(result_r[224*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001C2_AdderTree0000000001(.i_data({mult_result_i[224][3],mult_result_i[224][2],mult_result_i[224][1],mult_result_i[224][0]}), .o_data(result_i[224*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001C3_AdderTree0000000001(.i_data({mult_result_r[225][3],mult_result_r[225][2],mult_result_r[225][1],mult_result_r[225][0]}), .o_data(result_r[225*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001C4_AdderTree0000000001(.i_data({mult_result_i[225][3],mult_result_i[225][2],mult_result_i[225][1],mult_result_i[225][0]}), .o_data(result_i[225*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001C5_AdderTree0000000001(.i_data({mult_result_r[226][3],mult_result_r[226][2],mult_result_r[226][1],mult_result_r[226][0]}), .o_data(result_r[226*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001C6_AdderTree0000000001(.i_data({mult_result_i[226][3],mult_result_i[226][2],mult_result_i[226][1],mult_result_i[226][0]}), .o_data(result_i[226*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001C7_AdderTree0000000001(.i_data({mult_result_r[227][3],mult_result_r[227][2],mult_result_r[227][1],mult_result_r[227][0]}), .o_data(result_r[227*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001C8_AdderTree0000000001(.i_data({mult_result_i[227][3],mult_result_i[227][2],mult_result_i[227][1],mult_result_i[227][0]}), .o_data(result_i[227*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001C9_AdderTree0000000001(.i_data({mult_result_r[228][3],mult_result_r[228][2],mult_result_r[228][1],mult_result_r[228][0]}), .o_data(result_r[228*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001CA_AdderTree0000000001(.i_data({mult_result_i[228][3],mult_result_i[228][2],mult_result_i[228][1],mult_result_i[228][0]}), .o_data(result_i[228*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001CB_AdderTree0000000001(.i_data({mult_result_r[229][3],mult_result_r[229][2],mult_result_r[229][1],mult_result_r[229][0]}), .o_data(result_r[229*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001CC_AdderTree0000000001(.i_data({mult_result_i[229][3],mult_result_i[229][2],mult_result_i[229][1],mult_result_i[229][0]}), .o_data(result_i[229*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001CD_AdderTree0000000001(.i_data({mult_result_r[230][3],mult_result_r[230][2],mult_result_r[230][1],mult_result_r[230][0]}), .o_data(result_r[230*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001CE_AdderTree0000000001(.i_data({mult_result_i[230][3],mult_result_i[230][2],mult_result_i[230][1],mult_result_i[230][0]}), .o_data(result_i[230*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001CF_AdderTree0000000001(.i_data({mult_result_r[231][3],mult_result_r[231][2],mult_result_r[231][1],mult_result_r[231][0]}), .o_data(result_r[231*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001D0_AdderTree0000000001(.i_data({mult_result_i[231][3],mult_result_i[231][2],mult_result_i[231][1],mult_result_i[231][0]}), .o_data(result_i[231*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001D1_AdderTree0000000001(.i_data({mult_result_r[232][3],mult_result_r[232][2],mult_result_r[232][1],mult_result_r[232][0]}), .o_data(result_r[232*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001D2_AdderTree0000000001(.i_data({mult_result_i[232][3],mult_result_i[232][2],mult_result_i[232][1],mult_result_i[232][0]}), .o_data(result_i[232*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001D3_AdderTree0000000001(.i_data({mult_result_r[233][3],mult_result_r[233][2],mult_result_r[233][1],mult_result_r[233][0]}), .o_data(result_r[233*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001D4_AdderTree0000000001(.i_data({mult_result_i[233][3],mult_result_i[233][2],mult_result_i[233][1],mult_result_i[233][0]}), .o_data(result_i[233*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001D5_AdderTree0000000001(.i_data({mult_result_r[234][3],mult_result_r[234][2],mult_result_r[234][1],mult_result_r[234][0]}), .o_data(result_r[234*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001D6_AdderTree0000000001(.i_data({mult_result_i[234][3],mult_result_i[234][2],mult_result_i[234][1],mult_result_i[234][0]}), .o_data(result_i[234*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001D7_AdderTree0000000001(.i_data({mult_result_r[235][3],mult_result_r[235][2],mult_result_r[235][1],mult_result_r[235][0]}), .o_data(result_r[235*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001D8_AdderTree0000000001(.i_data({mult_result_i[235][3],mult_result_i[235][2],mult_result_i[235][1],mult_result_i[235][0]}), .o_data(result_i[235*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001D9_AdderTree0000000001(.i_data({mult_result_r[236][3],mult_result_r[236][2],mult_result_r[236][1],mult_result_r[236][0]}), .o_data(result_r[236*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001DA_AdderTree0000000001(.i_data({mult_result_i[236][3],mult_result_i[236][2],mult_result_i[236][1],mult_result_i[236][0]}), .o_data(result_i[236*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001DB_AdderTree0000000001(.i_data({mult_result_r[237][3],mult_result_r[237][2],mult_result_r[237][1],mult_result_r[237][0]}), .o_data(result_r[237*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001DC_AdderTree0000000001(.i_data({mult_result_i[237][3],mult_result_i[237][2],mult_result_i[237][1],mult_result_i[237][0]}), .o_data(result_i[237*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001DD_AdderTree0000000001(.i_data({mult_result_r[238][3],mult_result_r[238][2],mult_result_r[238][1],mult_result_r[238][0]}), .o_data(result_r[238*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001DE_AdderTree0000000001(.i_data({mult_result_i[238][3],mult_result_i[238][2],mult_result_i[238][1],mult_result_i[238][0]}), .o_data(result_i[238*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001DF_AdderTree0000000001(.i_data({mult_result_r[239][3],mult_result_r[239][2],mult_result_r[239][1],mult_result_r[239][0]}), .o_data(result_r[239*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001E0_AdderTree0000000001(.i_data({mult_result_i[239][3],mult_result_i[239][2],mult_result_i[239][1],mult_result_i[239][0]}), .o_data(result_i[239*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001E1_AdderTree0000000001(.i_data({mult_result_r[240][3],mult_result_r[240][2],mult_result_r[240][1],mult_result_r[240][0]}), .o_data(result_r[240*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001E2_AdderTree0000000001(.i_data({mult_result_i[240][3],mult_result_i[240][2],mult_result_i[240][1],mult_result_i[240][0]}), .o_data(result_i[240*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001E3_AdderTree0000000001(.i_data({mult_result_r[241][3],mult_result_r[241][2],mult_result_r[241][1],mult_result_r[241][0]}), .o_data(result_r[241*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001E4_AdderTree0000000001(.i_data({mult_result_i[241][3],mult_result_i[241][2],mult_result_i[241][1],mult_result_i[241][0]}), .o_data(result_i[241*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001E5_AdderTree0000000001(.i_data({mult_result_r[242][3],mult_result_r[242][2],mult_result_r[242][1],mult_result_r[242][0]}), .o_data(result_r[242*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001E6_AdderTree0000000001(.i_data({mult_result_i[242][3],mult_result_i[242][2],mult_result_i[242][1],mult_result_i[242][0]}), .o_data(result_i[242*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001E7_AdderTree0000000001(.i_data({mult_result_r[243][3],mult_result_r[243][2],mult_result_r[243][1],mult_result_r[243][0]}), .o_data(result_r[243*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001E8_AdderTree0000000001(.i_data({mult_result_i[243][3],mult_result_i[243][2],mult_result_i[243][1],mult_result_i[243][0]}), .o_data(result_i[243*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001E9_AdderTree0000000001(.i_data({mult_result_r[244][3],mult_result_r[244][2],mult_result_r[244][1],mult_result_r[244][0]}), .o_data(result_r[244*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001EA_AdderTree0000000001(.i_data({mult_result_i[244][3],mult_result_i[244][2],mult_result_i[244][1],mult_result_i[244][0]}), .o_data(result_i[244*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001EB_AdderTree0000000001(.i_data({mult_result_r[245][3],mult_result_r[245][2],mult_result_r[245][1],mult_result_r[245][0]}), .o_data(result_r[245*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001EC_AdderTree0000000001(.i_data({mult_result_i[245][3],mult_result_i[245][2],mult_result_i[245][1],mult_result_i[245][0]}), .o_data(result_i[245*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001ED_AdderTree0000000001(.i_data({mult_result_r[246][3],mult_result_r[246][2],mult_result_r[246][1],mult_result_r[246][0]}), .o_data(result_r[246*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001EE_AdderTree0000000001(.i_data({mult_result_i[246][3],mult_result_i[246][2],mult_result_i[246][1],mult_result_i[246][0]}), .o_data(result_i[246*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001EF_AdderTree0000000001(.i_data({mult_result_r[247][3],mult_result_r[247][2],mult_result_r[247][1],mult_result_r[247][0]}), .o_data(result_r[247*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001F0_AdderTree0000000001(.i_data({mult_result_i[247][3],mult_result_i[247][2],mult_result_i[247][1],mult_result_i[247][0]}), .o_data(result_i[247*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001F1_AdderTree0000000001(.i_data({mult_result_r[248][3],mult_result_r[248][2],mult_result_r[248][1],mult_result_r[248][0]}), .o_data(result_r[248*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001F2_AdderTree0000000001(.i_data({mult_result_i[248][3],mult_result_i[248][2],mult_result_i[248][1],mult_result_i[248][0]}), .o_data(result_i[248*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001F3_AdderTree0000000001(.i_data({mult_result_r[249][3],mult_result_r[249][2],mult_result_r[249][1],mult_result_r[249][0]}), .o_data(result_r[249*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001F4_AdderTree0000000001(.i_data({mult_result_i[249][3],mult_result_i[249][2],mult_result_i[249][1],mult_result_i[249][0]}), .o_data(result_i[249*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001F5_AdderTree0000000001(.i_data({mult_result_r[250][3],mult_result_r[250][2],mult_result_r[250][1],mult_result_r[250][0]}), .o_data(result_r[250*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001F6_AdderTree0000000001(.i_data({mult_result_i[250][3],mult_result_i[250][2],mult_result_i[250][1],mult_result_i[250][0]}), .o_data(result_i[250*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001F7_AdderTree0000000001(.i_data({mult_result_r[251][3],mult_result_r[251][2],mult_result_r[251][1],mult_result_r[251][0]}), .o_data(result_r[251*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001F8_AdderTree0000000001(.i_data({mult_result_i[251][3],mult_result_i[251][2],mult_result_i[251][1],mult_result_i[251][0]}), .o_data(result_i[251*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001F9_AdderTree0000000001(.i_data({mult_result_r[252][3],mult_result_r[252][2],mult_result_r[252][1],mult_result_r[252][0]}), .o_data(result_r[252*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001FA_AdderTree0000000001(.i_data({mult_result_i[252][3],mult_result_i[252][2],mult_result_i[252][1],mult_result_i[252][0]}), .o_data(result_i[252*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001FB_AdderTree0000000001(.i_data({mult_result_r[253][3],mult_result_r[253][2],mult_result_r[253][1],mult_result_r[253][0]}), .o_data(result_r[253*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001FC_AdderTree0000000001(.i_data({mult_result_i[253][3],mult_result_i[253][2],mult_result_i[253][1],mult_result_i[253][0]}), .o_data(result_i[253*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001FD_AdderTree0000000001(.i_data({mult_result_r[254][3],mult_result_r[254][2],mult_result_r[254][1],mult_result_r[254][0]}), .o_data(result_r[254*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001FE_AdderTree0000000001(.i_data({mult_result_i[254][3],mult_result_i[254][2],mult_result_i[254][1],mult_result_i[254][0]}), .o_data(result_i[254*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_00000001FF_AdderTree0000000001(.i_data({mult_result_r[255][3],mult_result_r[255][2],mult_result_r[255][1],mult_result_r[255][0]}), .o_data(result_r[255*12+:12]), .i_clk(i_clk));
AdderTree0000000001  u_0000000200_AdderTree0000000001(.i_data({mult_result_i[255][3],mult_result_i[255][2],mult_result_i[255][1],mult_result_i[255][0]}), .o_data(result_i[255*12+:12]), .i_clk(i_clk));
 endmodule
