 module Delay0000000004 (
    i_data, o_data
 );
 // Input and output ports
 input [13-1:0] i_data;
 output [13-1:0] o_data;
 assign o_data = i_data;
 endmodule
