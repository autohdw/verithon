 module TOP #(vparam_top1, vparam_top2, vparam_top3)(
 port_top1,
 port_top2,
 );
MUL #(.vparam1(3), .vparam2(6), .vparamN(5)) MUL1 (.PORT1(aaa), .PORT2(bbb), .PORT3(ccc));
 start of module TOP
 middle of module TOP
 end of module TOP
 endmodule
