 module Delay000000000A (
    i_data, o_data
 );
 // Input and output ports
 input [12-1:0] i_data;
 output [12-1:0] o_data;
 assign o_data = i_data;
 endmodule
