 module Delay000000000B (
    i_data, o_data
 );
 // Input and output ports
 input [16-1:0] i_data;
 output [16-1:0] o_data;
 assign o_data = i_data;
 endmodule
